
/* Source file "
	partitionlib/uvm_custom_install_verdi_recording_zILyrc/uvm_custom_install_verdi_recording.v
	", line 1 */
(* VCS_LogicalLibrary = "VCS_PARTCOMP_LIB" *)
config pc_uvm_custom_install_verdi_recording_config;
	design pc_uvm_custom_install_verdi_recording DEFAULT.
		uvm_custom_install_verdi_recording DEFAULT.Risc_16_bit_test;
	cell uvm_custom_install_verdi_recording liblist DEFAULT;
	cell Risc_16_bit_test liblist DEFAULT;
	instance Risc_16_bit_test.dut use VCS_PARTCOMP_LIB.Risc_16_bit_g2J7Bb;
	partition instance Risc_16_bit_test.dut;
endconfig
`timescale 1ns/1fs
/* Source file "", line 0 */

(* PARTCOMP_WRAPPER = 1, PARTCOMP_DOLLAR_UNIT = "DEFAULT._vcs_unit__17393910" *)

(* VCS_LogicalLibrary = "VCS_PARTCOMP_LIB" *)

`timescale 1ns/1fs
(* orig_name = "pc_uvm_custom_install_verdi_recording" *)
module pc_uvm_custom_install_verdi_recording;


	wire			__vcs_0_SI_DT6vKb;
	wire			__vcs_1_SI_DT6vKb;
	wire			__vcs_2_SI_DT6vKb;
	wire			__vcs_3_SI_DT6vKb;
	wire			__vcs_4_SI_DT6vKb;
	wire			__vcs_5_SI_DT6vKb;
	wire			__vcs_6_SI_DT6vKb;
	wire			__vcs_7_SI_DT6vKb;
	wire			__vcs_8_SI_DT6vKb;
	wire			__vcs_9_SI_DT6vKb;
	wire			__vcs_A_QN_DT6vKb;
	wire			__vcs_B_SI_DT6vKb;
	wire			__vcs_C_SI_DT6vKb;
	wire			__vcs_D_SI_DT6vKb;
	wire			__vcs_E_SI_DT6vKb;
	wire			__vcs_F_SI_DT6vKb;
	wire			__vcs_10_SI_DT6vKb;
	wire			__vcs_11_SI_DT6vKb;
	wire			__vcs_12_Q_DT6vKb;
	wire			__vcs_13_QN_DT6vKb;
	wire			__vcs_14_QN_DT6vKb;
	wire			__vcs_15_QN_DT6vKb;
	wire			__vcs_16_QN_DT6vKb;
	wire			__vcs_17_QN_DT6vKb;
	wire			__vcs_18_QN_DT6vKb;
	wire			__vcs_19_QN_DT6vKb;
	wire			__vcs_1A_QN_DT6vKb;
	wire			__vcs_1B_QN_DT6vKb;
	wire			__vcs_1C_QN_DT6vKb;
	wire			__vcs_1D_QN_DT6vKb;
	wire			__vcs_1E_QN_DT6vKb;
	wire			__vcs_1F_QN_DT6vKb;
	wire			__vcs_20_QN_DT6vKb;
	wire			__vcs_21_QN_DT6vKb;
	wire			__vcs_22_QN_DT6vKb;
	wire			__vcs_23_QN_DT6vKb;
	wire			__vcs_24_SI_DT6vKb;
	wire			__vcs_25_QN_DT6vKb;
	wire			__vcs_26_Q_DT6vKb;
	wire			__vcs_27_QN_DT6vKb;
	wire			__vcs_28_Q_DT6vKb;
	wire			__vcs_29_SI_DT6vKb;
	wire			__vcs_2A_SI_DT6vKb;
	wire			__vcs_2B_Q_DT6vKb;
	wire			__vcs_2C_SI_DT6vKb;
	wire			__vcs_2D_QN_DT6vKb;
	wire			__vcs_2E_SI_DT6vKb;
	wire			__vcs_2F_QN_DT6vKb;
	wire			__vcs_30_QN_DT6vKb;
	wire			__vcs_31_SI_DT6vKb;
	wire			__vcs_32_QN_DT6vKb;
	wire			__vcs_33_SI_DT6vKb;
	wire			__vcs_34_SI_DT6vKb;
	wire			__vcs_35_SI_DT6vKb;
	wire			__vcs_36_SI_DT6vKb;
	wire			__vcs_37_SI_DT6vKb;
	wire			__vcs_38_SI_DT6vKb;
	wire			__vcs_39_SI_DT6vKb;
	wire			__vcs_3A_SI_DT6vKb;
	wire			__vcs_3B_SI_DT6vKb;
	wire			__vcs_3C_SI_DT6vKb;
	wire			__vcs_3D_SI_DT6vKb;
	wire			__vcs_3E_SI_DT6vKb;
	wire			__vcs_3F_SI_DT6vKb;
	wire			__vcs_40_SI_DT6vKb;
	wire			__vcs_41_SI_DT6vKb;
	wire			__vcs_42_QN_DT6vKb;
	wire			__vcs_43_SI_DT6vKb;
	wire			__vcs_44_SI_DT6vKb;
	wire			__vcs_45_SI_DT6vKb;
	wire			__vcs_46_SI_DT6vKb;
	wire			__vcs_47_SI_DT6vKb;
	wire			__vcs_48_QN_DT6vKb;
	wire			__vcs_49_QN_DT6vKb;
	wire			__vcs_4A_QN_DT6vKb;
	wire			__vcs_4B_QN_DT6vKb;
	wire			__vcs_4C_QN_DT6vKb;
	wire			__vcs_4D_QN_DT6vKb;
	wire			__vcs_4E_QN_DT6vKb;
	wire			__vcs_4F_QN_DT6vKb;
	wire			__vcs_50_QN_DT6vKb;
	wire			__vcs_51_QN_DT6vKb;
	wire			__vcs_52_SI_DT6vKb;
	wire			__vcs_53_SI_DT6vKb;
	wire			__vcs_54_SI_DT6vKb;
	wire			__vcs_55_SI_DT6vKb;
	wire			__vcs_56_QN_DT6vKb;
	wire			__vcs_57_QN_DT6vKb;
	wire			__vcs_58_QN_DT6vKb;
	wire			__vcs_59_SI_DT6vKb;
	wire			__vcs_5A_SI_DT6vKb;
	wire			__vcs_5B_SI_DT6vKb;
	wire			__vcs_5C_SI_DT6vKb;
	wire			__vcs_5D_SI_DT6vKb;
	wire			__vcs_5E_SI_DT6vKb;
	wire			__vcs_5F_SI_DT6vKb;
	wire			__vcs_60_SI_DT6vKb;
	wire			__vcs_61_SI_DT6vKb;
	wire			__vcs_62_SI_DT6vKb;
	wire			__vcs_63_SI_DT6vKb;
	wire			__vcs_64_QN_DT6vKb;
	wire			__vcs_65_SI_DT6vKb;
	wire			__vcs_66_QN_DT6vKb;
	wire			__vcs_67_QN_DT6vKb;
	wire			__vcs_68_QN_DT6vKb;
	wire			__vcs_69_QN_DT6vKb;
	wire			__vcs_6A_QN_DT6vKb;
	wire			__vcs_6B_QN_DT6vKb;
	wire			__vcs_6C_QN_DT6vKb;
	wire			__vcs_6D_QN_DT6vKb;
	wire			__vcs_6E_QN_DT6vKb;
	wire			__vcs_6F_SI_DT6vKb;
	wire			__vcs_70_SI_DT6vKb;
	wire			__vcs_71_SI_DT6vKb;
	wire			__vcs_72_D_DT6vKb;
	wire			__vcs_73_QN_DT6vKb;
	wire			__vcs_74_SI_DT6vKb;
	wire			__vcs_75_SI_DT6vKb;
	wire			__vcs_76_SI_DT6vKb;
	wire			__vcs_77_SI_DT6vKb;
	wire			__vcs_78_SI_DT6vKb;
	wire			__vcs_79_Q_DT6vKb;
	wire			__vcs_7A_SI_DT6vKb;
	wire			__vcs_7B_SI_DT6vKb;
	wire			__vcs_7C_SI_DT6vKb;
	wire			__vcs_7D_SI_DT6vKb;
	wire			__vcs_7E_D_DT6vKb;
	wire			__vcs_7F_QN_DT6vKb;
	wire			__vcs_80_SI_DT6vKb;
	wire			__vcs_81_SI_DT6vKb;
	wire			__vcs_82_QN_DT6vKb;
	wire			__vcs_83_QN_DT6vKb;
	wire			__vcs_84_QN_DT6vKb;
	wire			__vcs_85_QN_DT6vKb;
	wire			__vcs_86_QN_DT6vKb;
	wire			__vcs_87_QN_DT6vKb;
	wire			__vcs_88_QN_DT6vKb;
	wire			__vcs_89_QN_DT6vKb;
	wire			__vcs_8A_SI_DT6vKb;
	wire			__vcs_8B_Q_DT6vKb;
	wire			__vcs_8C_D_DT6vKb;
	wire			__vcs_8D_Q_DT6vKb;
	wire			__vcs_8E_SI_DT6vKb;
	wire			__vcs_8F_Q_DT6vKb;
	wire			__vcs_90_Q_DT6vKb;
	wire			__vcs_91_SI_DT6vKb;
	wire			__vcs_92_Q_DT6vKb;
	wire			__vcs_93_D_DT6vKb;
	wire			__vcs_94_SI_DT6vKb;
	wire			__vcs_95_SI_DT6vKb;
	wire			__vcs_96_SI_DT6vKb;
	wire			__vcs_97_SI_DT6vKb;
	wire			__vcs_98_SI_DT6vKb;
	wire			__vcs_99_SI_DT6vKb;
	wire			__vcs_9A_SI_DT6vKb;
	wire			__vcs_9B_SI_DT6vKb;
	wire			__vcs_9C_Q_DT6vKb;
	wire			__vcs_9D_QN_DT6vKb;
	wire			__vcs_9E_QN_DT6vKb;
	wire			__vcs_9F_QN_DT6vKb;
	wire			__vcs_A0_QN_DT6vKb;
	wire			__vcs_A1_Q_DT6vKb;
	wire			__vcs_A2_QN_DT6vKb;
	wire			__vcs_A3_QN_DT6vKb;
	wire			__vcs_A4_QN_DT6vKb;
	wire			__vcs_A5_QN_DT6vKb;
	wire			__vcs_A6_QN_DT6vKb;
	wire			__vcs_A7_SI_DT6vKb;
	wire			__vcs_A8_SI_DT6vKb;
	wire			__vcs_A9_SI_DT6vKb;
	wire			__vcs_AA_SI_DT6vKb;
	wire			__vcs_AB_SI_DT6vKb;
	wire			__vcs_AC_SI_DT6vKb;
	wire			__vcs_AD_SI_DT6vKb;
	wire			__vcs_AE_SI_DT6vKb;
	wire			__vcs_AF_SI_DT6vKb;
	wire			__vcs_B0_QN_DT6vKb;
	wire			__vcs_B1_QN_DT6vKb;
	wire			__vcs_B2_QN_DT6vKb;
	wire			__vcs_B3_QN_DT6vKb;
	wire			__vcs_B4_QN_DT6vKb;
	wire			__vcs_B5_QN_DT6vKb;
	wire			__vcs_B6_QN_DT6vKb;
	wire			__vcs_B7_QN_DT6vKb;
	wire			__vcs_B8_QN_DT6vKb;
	wire			__vcs_B9_SI_DT6vKb;
	wire			__vcs_BA_QN_DT6vKb;
	wire			__vcs_BB_QN_DT6vKb;
	wire			__vcs_BC_SI_DT6vKb;
	wire			__vcs_BD_SI_DT6vKb;
	wire			__vcs_BE_SI_DT6vKb;
	wire			__vcs_BF_SI_DT6vKb;
	wire			__vcs_C0_SI_DT6vKb;
	wire			__vcs_C1_QN_DT6vKb;
	wire			__vcs_C2_SI_DT6vKb;
	wire			__vcs_C3_SI_DT6vKb;
	wire			__vcs_C4_SI_DT6vKb;
	wire			__vcs_C5_SI_DT6vKb;
	wire			__vcs_C6_QN_DT6vKb;
	wire			__vcs_C7_SI_DT6vKb;
	wire			__vcs_C8_QN_DT6vKb;
	wire			__vcs_C9_QN_DT6vKb;
	wire			__vcs_CA_QN_DT6vKb;
	wire			__vcs_CB_QN_DT6vKb;
	wire			__vcs_CC_QN_DT6vKb;
	wire			__vcs_CD_SI_DT6vKb;
	wire			__vcs_CE_QN_DT6vKb;
	wire			__vcs_CF_QN_DT6vKb;
	wire			__vcs_D0_QN_DT6vKb;
	wire			__vcs_D1_SI_DT6vKb;
	wire			__vcs_D2_QN_DT6vKb;
	wire			__vcs_D3_QN_DT6vKb;
	wire			__vcs_D4_QN_DT6vKb;
	wire			__vcs_D5_SI_DT6vKb;
	wire			__vcs_D6_SI_DT6vKb;
	wire			__vcs_D7_QN_DT6vKb;
	wire			__vcs_D8_SI_DT6vKb;
	wire			__vcs_D9_SI_DT6vKb;
	wire			__vcs_DA_Q_DT6vKb;
	wire			__vcs_DB_SI_DT6vKb;
	wire			__vcs_DC_SI_DT6vKb;
	wire			__vcs_DD_SI_DT6vKb;
	wire			__vcs_DE_QN_DT6vKb;
	wire			__vcs_DF_SI_DT6vKb;
	wire			__vcs_E0_SI_DT6vKb;
	wire			__vcs_E1_SI_DT6vKb;
	wire			__vcs_E2_QN_DT6vKb;
	wire			__vcs_E3_SI_DT6vKb;
	wire			__vcs_E4_Q_DT6vKb;
	wire			__vcs_E5_QN_DT6vKb;
	wire			__vcs_E6_Q_DT6vKb;
	wire			__vcs_E7_SI_DT6vKb;
	wire			__vcs_E8_QN_DT6vKb;
	wire			__vcs_E9_QN_DT6vKb;
	wire			__vcs_EA_QN_DT6vKb;
	wire			__vcs_EB_QN_DT6vKb;
	wire			__vcs_EC_QN_DT6vKb;
	wire			__vcs_ED_SI_DT6vKb;
	wire			__vcs_EE_QN_DT6vKb;
	wire			__vcs_EF_QN_DT6vKb;
	wire			__vcs_F0_QN_DT6vKb;
	wire			__vcs_F1_QN_DT6vKb;
	wire			__vcs_F2_SI_DT6vKb;
	wire			__vcs_F3_Q_DT6vKb;
	wire			__vcs_F4_QN_DT6vKb;
	wire			__vcs_F5_QN_DT6vKb;
	wire			__vcs_F6_SI_DT6vKb;
	wire			__vcs_F7_QN_DT6vKb;
	wire			__vcs_F8_SI_DT6vKb;
	wire			__vcs_F9_SI_DT6vKb;
	wire			__vcs_FA_QN_DT6vKb;
	wire			__vcs_FB_SI_DT6vKb;
	wire			__vcs_FC_SI_DT6vKb;
	wire			__vcs_FD_SI_DT6vKb;
	wire			__vcs_FE_SI_DT6vKb;
	wire			__vcs_FF_SI_DT6vKb;
	wire			__vcs_100_QN_DT6vKb;
	wire			__vcs_101_SI_DT6vKb;
	wire			__vcs_102_SI_DT6vKb;
	wire			__vcs_103_SI_DT6vKb;
	wire			__vcs_104_SI_DT6vKb;
	wire			__vcs_105_SI_DT6vKb;
	wire			__vcs_106_QN_DT6vKb;
	wire			__vcs_107_QN_DT6vKb;
	wire			__vcs_108_SI_DT6vKb;
	wire			__vcs_109_QN_DT6vKb;
	wire			__vcs_10A_QN_DT6vKb;
	wire			__vcs_10B_QN_DT6vKb;
	wire			__vcs_10C_QN_DT6vKb;
	wire			__vcs_10D_QN_DT6vKb;
	wire			__vcs_10E_QN_DT6vKb;
	wire			__vcs_10F_SI_DT6vKb;
	wire			__vcs_110_QN_DT6vKb;
	wire			__vcs_111_QN_DT6vKb;
	wire			__vcs_112_QN_DT6vKb;
	wire			__vcs_113_QN_DT6vKb;
	wire			__vcs_114_SI_DT6vKb;
	wire			__vcs_115_QN_DT6vKb;
	wire			__vcs_116_QN_DT6vKb;
	wire			__vcs_117_SI_DT6vKb;
	wire			__vcs_118_QN_DT6vKb;
	wire			__vcs_119_SI_DT6vKb;
	wire			__vcs_11A_SI_DT6vKb;
	wire			__vcs_11B_QN_DT6vKb;
	wire			__vcs_11C_SI_DT6vKb;
	wire			__vcs_11D_SI_DT6vKb;
	wire			__vcs_11E_SI_DT6vKb;
	wire			__vcs_11F_SI_DT6vKb;
	wire			__vcs_120_SI_DT6vKb;
	wire			__vcs_121_QN_DT6vKb;
	wire			__vcs_122_SI_DT6vKb;
	wire			__vcs_123_SI_DT6vKb;
	wire			__vcs_124_SI_DT6vKb;
	wire			__vcs_125_SI_DT6vKb;
	wire			__vcs_126_SI_DT6vKb;
	wire			__vcs_127_QN_DT6vKb;
	wire			__vcs_128_QN_DT6vKb;
	wire			__vcs_129_SI_DT6vKb;
	wire			__vcs_12A_QN_DT6vKb;
	wire			__vcs_12B_QN_DT6vKb;
	wire			__vcs_12C_QN_DT6vKb;
	wire			__vcs_12D_QN_DT6vKb;
	wire			__vcs_12E_QN_DT6vKb;
	wire			__vcs_12F_SI_DT6vKb;
	wire			__vcs_130_QN_DT6vKb;
	wire			__vcs_131_QN_DT6vKb;
	wire			__vcs_132_QN_DT6vKb;
	wire			__vcs_133_QN_DT6vKb;
	wire			__vcs_134_QN_DT6vKb;
	wire			__vcs_135_QN_DT6vKb;
	wire			__vcs_136_QN_DT6vKb;
	wire			__vcs_137_QN_DT6vKb;
	wire			__vcs_138_SI_DT6vKb;
	wire			__vcs_139_QN_DT6vKb;
	wire			__vcs_13A_QN_DT6vKb;
	wire			__vcs_13B_QN_DT6vKb;
	wire			__vcs_13C_QN_DT6vKb;
	wire			__vcs_13D_QN_DT6vKb;
	wire			__vcs_13E_QN_DT6vKb;
	wire			__vcs_13F_SI_DT6vKb;
	wire			__vcs_140_QN_DT6vKb;
	wire			__vcs_141_QN_DT6vKb;
	wire			__vcs_142_SI_DT6vKb;
	wire			__vcs_143_QN_DT6vKb;
	wire			__vcs_144_SI_DT6vKb;
	wire			__vcs_145_SI_DT6vKb;
	wire			__vcs_146_QN_DT6vKb;
	wire			__vcs_147_SI_DT6vKb;
	wire			__vcs_148_SI_DT6vKb;
	wire			__vcs_149_QN_DT6vKb;
	wire			__vcs_14A_SI_DT6vKb;
	wire			__vcs_14B_SI_DT6vKb;
	wire			__vcs_14C_SI_DT6vKb;
	wire			__vcs_14D_SI_DT6vKb;
	wire			__vcs_14E_SI_DT6vKb;
	wire			__vcs_14F_SI_DT6vKb;
	wire			__vcs_150_SI_DT6vKb;
	wire			__vcs_151_SI_DT6vKb;
	wire			__vcs_152_SI_DT6vKb;
	wire			__vcs_153_SI_DT6vKb;
	wire			__vcs_154_SI_DT6vKb;
	wire			__vcs_155_QN_DT6vKb;
	wire			__vcs_156_SI_DT6vKb;
	wire			__vcs_157_SI_DT6vKb;
	wire			__vcs_158_SI_DT6vKb;
	wire			__vcs_159_SI_DT6vKb;
	wire			__vcs_15A_SI_DT6vKb;
	wire			__vcs_15B_SI_DT6vKb;
	wire			__vcs_15C_QN_DT6vKb;
	wire			__vcs_15D_QN_DT6vKb;
	wire			__vcs_15E_SI_DT6vKb;
	wire			__vcs_15F_SI_DT6vKb;
	wire			__vcs_160_QN_DT6vKb;
	wire			__vcs_161_QN_DT6vKb;
	wire			__vcs_162_QN_DT6vKb;
	wire			__vcs_163_SI_DT6vKb;
	wire			__vcs_164_QN_DT6vKb;
	wire			__vcs_165_QN_DT6vKb;
	wire			__vcs_166_QN_DT6vKb;
	wire			__vcs_167_QN_DT6vKb;
	wire			__vcs_168_QN_DT6vKb;
	wire			__vcs_169_QN_DT6vKb;
	wire			__vcs_16A_QN_DT6vKb;
	wire			__vcs_16B_QN_DT6vKb;
	wire			__vcs_16C_QN_DT6vKb;
	wire			__vcs_16D_QN_DT6vKb;
	wire			__vcs_16E_SI_DT6vKb;
	wire			__vcs_16F_QN_DT6vKb;
	wire			__vcs_170_QN_DT6vKb;
	wire			__vcs_171_QN_DT6vKb;
	wire			__vcs_172_QN_DT6vKb;
	wire			__vcs_173_QN_DT6vKb;
	wire			__vcs_174_SI_DT6vKb;
	wire			__vcs_175_QN_DT6vKb;
	wire			__vcs_176_QN_DT6vKb;
	wire			__vcs_177_SI_DT6vKb;
	wire			__vcs_178_SI_DT6vKb;
	wire			__vcs_179_Q_DT6vKb;
	wire			__vcs_17A_SI_DT6vKb;
	wire			__vcs_17B_QN_DT6vKb;
	wire			__vcs_17C_QN_DT6vKb;
	wire			__vcs_17D_SI_DT6vKb;
	wire			__vcs_17E_QN_DT6vKb;
	wire			__vcs_17F_SI_DT6vKb;
	wire			__vcs_180_SI_DT6vKb;
	wire			__vcs_181_SI_DT6vKb;
	wire			__vcs_182_QN_DT6vKb;
	wire			__vcs_183_Q_DT6vKb;
	wire			__vcs_184_SI_DT6vKb;
	wire			__vcs_185_SI_DT6vKb;
	wire			__vcs_186_SI_DT6vKb;
	wire			__vcs_187_SI_DT6vKb;
	wire			__vcs_188_SI_DT6vKb;
	wire			__vcs_189_SI_DT6vKb;
	wire			__vcs_18A_SI_DT6vKb;
	wire			__vcs_18B_SI_DT6vKb;
	wire			__vcs_18C_QN_DT6vKb;
	wire			__vcs_18D_SI_DT6vKb;
	wire			__vcs_18E_SI_DT6vKb;
	wire			__vcs_18F_SI_DT6vKb;
	wire			__vcs_190_SI_DT6vKb;
	wire			__vcs_191_SI_DT6vKb;
	wire			__vcs_192_SI_DT6vKb;
	wire			__vcs_193_SI_DT6vKb;
	wire			__vcs_194_SI_DT6vKb;
	wire			__vcs_195_SI_DT6vKb;
	wire			__vcs_196_QN_DT6vKb;
	wire			__vcs_197_SI_DT6vKb;
	wire			__vcs_198_QN_DT6vKb;
	wire			__vcs_199_QN_DT6vKb;
	wire			__vcs_19A_QN_DT6vKb;
	wire			__vcs_19B_QN_DT6vKb;
	wire			__vcs_19C_QN_DT6vKb;
	wire			__vcs_19D_QN_DT6vKb;
	wire			__vcs_19E_SI_DT6vKb;
	wire			__vcs_19F_QN_DT6vKb;
	wire			__vcs_1A0_QN_DT6vKb;
	wire			__vcs_1A1_QN_DT6vKb;
	wire			__vcs_1A2_QN_DT6vKb;
	wire			__vcs_1A3_QN_DT6vKb;
	wire			__vcs_1A4_QN_DT6vKb;
	wire			__vcs_1A5_QN_DT6vKb;
	wire			__vcs_1A6_QN_DT6vKb;
	wire			__vcs_1A7_SI_DT6vKb;
	wire			__vcs_1A8_QN_DT6vKb;
	wire			__vcs_1A9_QN_DT6vKb;
	wire			__vcs_1AA_QN_DT6vKb;
	wire			__vcs_1AB_QN_DT6vKb;
	wire			__vcs_1AC_QN_DT6vKb;
	wire			__vcs_1AD_QN_DT6vKb;
	wire			__vcs_1AE_SI_DT6vKb;
	wire			__vcs_1AF_QN_DT6vKb;
	wire			__vcs_1B0_SI_DT6vKb;
	wire			__vcs_1B1_SI_DT6vKb;
	wire			__vcs_1B2_QN_DT6vKb;
	wire			__vcs_1B3_SI_DT6vKb;
	wire			__vcs_1B4_SI_DT6vKb;
	wire			__vcs_1B5_QN_DT6vKb;
	wire			__vcs_1B6_QN_DT6vKb;
	wire			__vcs_1B7_SI_DT6vKb;
	wire			__vcs_1B8_QN_DT6vKb;
	wire			__vcs_1B9_SI_DT6vKb;
	wire			__vcs_1BA_SI_DT6vKb;
	wire			__vcs_1BB_QN_DT6vKb;
	wire			__vcs_1BC_SI_DT6vKb;
	wire			__vcs_1BD_SI_DT6vKb;
	wire			__vcs_1BE_SI_DT6vKb;
	wire			__vcs_1BF_SI_DT6vKb;
	wire			__vcs_1C0_SI_DT6vKb;
	wire			__vcs_1C1_SI_DT6vKb;
	wire			__vcs_1C2_SI_DT6vKb;
	wire			__vcs_1C3_SI_DT6vKb;
	wire			__vcs_1C4_SI_DT6vKb;
	wire			__vcs_1C5_SI_DT6vKb;
	wire			__vcs_1C6_SI_DT6vKb;
	wire			__vcs_1C7_QN_DT6vKb;
	wire			__vcs_1C8_SI_DT6vKb;
	wire			__vcs_1C9_SI_DT6vKb;
	wire			__vcs_1CA_SI_DT6vKb;
	wire			__vcs_1CB_SI_DT6vKb;
	wire			__vcs_1CC_SI_DT6vKb;
	wire			__vcs_1CD_SI_DT6vKb;
	wire			__vcs_1CE_SI_DT6vKb;
	wire			__vcs_1CF_SI_DT6vKb;
	wire			__vcs_1D0_QN_DT6vKb;
	wire			__vcs_1D1_QN_DT6vKb;
	wire			__vcs_1D2_QN_DT6vKb;
	wire			__vcs_1D3_QN_DT6vKb;
	wire			__vcs_1D4_QN_DT6vKb;
	wire			__vcs_1D5_SI_DT6vKb;
	wire			__vcs_1D6_QN_DT6vKb;
	wire			__vcs_1D7_QN_DT6vKb;
	wire			__vcs_1D8_QN_DT6vKb;
	wire			__vcs_1D9_QN_DT6vKb;
	wire			__vcs_1DA_QN_DT6vKb;
	wire			__vcs_1DB_QN_DT6vKb;
	wire			__vcs_1DC_QN_DT6vKb;
	wire			__vcs_1DD_QN_DT6vKb;
	wire			__vcs_1DE_QN_DT6vKb;
	wire			__vcs_1DF_QN_DT6vKb;
	wire			__vcs_1E0_QN_DT6vKb;
	wire			__vcs_1E1_SI_DT6vKb;
	wire			__vcs_1E2_QN_DT6vKb;
	wire			__vcs_1E3_QN_DT6vKb;
	wire			__vcs_1E4_QN_DT6vKb;
	wire			__vcs_1E5_QN_DT6vKb;
	wire			__vcs_1E6_SI_DT6vKb;
	wire			__vcs_1E7_SI_DT6vKb;
	wire			__vcs_1E8_SI_DT6vKb;
	wire			__vcs_1E9_QN_DT6vKb;
	wire			__vcs_1EA_SI_DT6vKb;
	wire			__vcs_1EB_SI_DT6vKb;
	wire			__vcs_1EC_QN_DT6vKb;
	wire			__vcs_1ED_QN_DT6vKb;
	wire			__vcs_1EE_SI_DT6vKb;
	wire			__vcs_1EF_QN_DT6vKb;
	wire			__vcs_1F0_SI_DT6vKb;
	wire			__vcs_1F1_SI_DT6vKb;
	wire			__vcs_1F2_SI_DT6vKb;
	wire			__vcs_1F3_SI_DT6vKb;
	wire			__vcs_1F4_SI_DT6vKb;
	wire			__vcs_1F5_SI_DT6vKb;
	wire			__vcs_1F6_SI_DT6vKb;
	wire			__vcs_1F7_SI_DT6vKb;
	wire			__vcs_1F8_SI_DT6vKb;
	wire			__vcs_1F9_SI_DT6vKb;
	wire			__vcs_1FA_SI_DT6vKb;
	wire			__vcs_1FB_SI_DT6vKb;
	wire			__vcs_1FC_SI_DT6vKb;
	wire			__vcs_1FD_SI_DT6vKb;
	wire			__vcs_1FE_QN_DT6vKb;
	wire			__vcs_1FF_SI_DT6vKb;
	wire			__vcs_200_SI_DT6vKb;
	wire			__vcs_201_SI_DT6vKb;
	wire			__vcs_202_SI_DT6vKb;
	wire			__vcs_203_SI_DT6vKb;
	wire			__vcs_204_SI_DT6vKb;
	wire			__vcs_205_SI_DT6vKb;
	wire			__vcs_206_QN_DT6vKb;
	wire			__vcs_207_QN_DT6vKb;
	wire			__vcs_208_QN_DT6vKb;
	wire			__vcs_209_QN_DT6vKb;
	wire			__vcs_20A_QN_DT6vKb;
	wire			__vcs_20B_QN_DT6vKb;
	wire			__vcs_20C_QN_DT6vKb;
	wire			__vcs_20D_QN_DT6vKb;
	wire			__vcs_20E_QN_DT6vKb;
	wire			__vcs_20F_QN_DT6vKb;
	wire			__vcs_210_QN_DT6vKb;
	wire			__vcs_211_QN_DT6vKb;
	wire			__vcs_212_Q_DT6vKb;
	wire			__vcs_213_QN_DT6vKb;
	wire			__vcs_214_QN_DT6vKb;
	wire			__vcs_215_QN_DT6vKb;
	wire			__vcs_216_QN_DT6vKb;
	wire			__vcs_217_QN_DT6vKb;
	wire			__vcs_218_SI_DT6vKb;
	wire			__vcs_219_QN_DT6vKb;
	wire			__vcs_21A_QN_DT6vKb;
	wire			__vcs_21B_SI_DT6vKb;
	wire			__vcs_21C_SI_DT6vKb;
	wire			__vcs_21D_SI_DT6vKb;
	wire			__vcs_21E_QN_DT6vKb;
	wire			__vcs_21F_SI_DT6vKb;
	wire			__vcs_220_QN_DT6vKb;
	wire			__vcs_221_QN_DT6vKb;
	wire			__vcs_222_SI_DT6vKb;
	wire			__vcs_223_QN_DT6vKb;
	wire			__vcs_224_SI_DT6vKb;
	wire			__vcs_225_Q_DT6vKb;
	wire			__vcs_226_SI_DT6vKb;
	wire			__vcs_227_SI_DT6vKb;

	initial begin : XmrProcess
	  $$xmr_map_rel(0, "Risc_16_bit_test", __vcs_0_SI_DT6vKb, 
		  "dut.DU.dm.\\memory_reg[0][8] .SI", 4, __vcs_1_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][4] .SI", 4, 
		  __vcs_2_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][8] .SI", 4, 
		  __vcs_3_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][4] .SI", 4, 
		  __vcs_4_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][8] .SI", 4, 
		  __vcs_5_SI_DT6vKb, "dut.DU.\\pc_current_reg[5] .SI", 3, 
		  __vcs_6_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][4] .SI", 4, 
		  __vcs_7_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][8] .SI", 4, 
		  __vcs_8_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][13] .SI", 4, 
		  __vcs_9_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][4] .SI", 4, 
		  __vcs_A_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][12] .QN", 4, 
		  __vcs_B_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][8] .SI", 4, 
		  __vcs_C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][4] .SI", 4, 
		  __vcs_D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][8] .SI", 4, 
		  __vcs_E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][4] .SI", 4, 
		  __vcs_F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][8] .SI", 4, 
		  __vcs_10_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][14] .SI", 4, 
		  __vcs_11_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][8] .SI", 4, 
		  __vcs_12_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][5] .Q",
		  4, __vcs_13_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][5] .QN", 4, 
		  __vcs_14_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][13] .QN", 4, 
		  __vcs_15_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][9] .QN", 4, 
		  __vcs_16_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][5] .QN", 4, 
		  __vcs_17_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][9] .QN", 4, 
		  __vcs_18_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][5] .QN", 4, 
		  __vcs_19_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][9] .QN", 4, 
		  __vcs_1A_QN_DT6vKb, "dut.DU.\\pc_current_reg[6] .QN", 3, 
		  __vcs_1B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][5] .QN", 4, 
		  __vcs_1C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][9] .QN", 4, 
		  __vcs_1D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][14] .QN", 4, 
		  __vcs_1E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][5] .QN", 4, 
		  __vcs_1F_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][9] .QN", 4, 
		  __vcs_20_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][5] .QN", 4, 
		  __vcs_21_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][9] .QN", 4, 
		  __vcs_22_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][5] .QN", 4, 
		  __vcs_23_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][9] .QN", 4, 
		  __vcs_24_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][12] .SI", 4, 
		  __vcs_25_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][9] .QN", 4, 
		  __vcs_26_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][12] .Q", 4, 
		  __vcs_27_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][15] .QN", 4, 
		  __vcs_28_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][9] .Q",
		  4, __vcs_29_SI_DT6vKb, "dut.DU.\\pc_current_reg[13] .SI", 3, 
		  __vcs_2A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][13] .SI", 4, 
		  __vcs_2B_Q_DT6vKb, "dut.DU.dm.\\memory_reg[1][1] .Q", 4, 
		  __vcs_2C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][14] .SI", 4, 
		  __vcs_2D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][13] .QN", 4, 
		  __vcs_2E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][15] .SI", 4, 
		  __vcs_2F_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][14] .QN", 4, 
		  __vcs_30_QN_DT6vKb, "dut.DU.\\pc_current_reg[14] .QN", 3, 
		  __vcs_31_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][12] .SI", 4, 
		  __vcs_32_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][15] .QN", 4, 
		  __vcs_33_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][5] .SI", 4, 
		  __vcs_34_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][5] .SI", 4, 
		  __vcs_35_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][13] .SI", 4, 
		  __vcs_36_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][9] .SI", 4, 
		  __vcs_37_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][5] .SI", 4, 
		  __vcs_38_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][9] .SI", 4, 
		  __vcs_39_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][5] .SI", 4, 
		  __vcs_3A_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][9] .SI", 4, 
		  __vcs_3B_SI_DT6vKb, "dut.DU.\\pc_current_reg[6] .SI", 3, 
		  __vcs_3C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][5] .SI", 4, 
		  __vcs_3D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][9] .SI", 4, 
		  __vcs_3E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][14] .SI", 4, 
		  __vcs_3F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][5] .SI", 4, 
		  __vcs_40_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][9] .SI", 4, 
		  __vcs_41_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][5] .SI", 4, 
		  __vcs_42_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][13] .QN", 4, 
		  __vcs_43_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][9] .SI", 4, 
		  __vcs_44_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][5] .SI", 4, 
		  __vcs_45_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][9] .SI", 4, 
		  __vcs_46_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][9] .SI", 4, 
		  __vcs_47_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][15] .SI", 4, 
		  __vcs_48_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][14] .QN", 4, 
		  __vcs_49_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][6] .QN", 4, 
		  __vcs_4A_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][6] .QN", 4, 
		  __vcs_4B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][6] .QN", 4, 
		  __vcs_4C_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][6] .QN", 4, 
		  __vcs_4D_QN_DT6vKb, "dut.DU.\\pc_current_reg[7] .QN", 3, 
		  __vcs_4E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][6] .QN", 4, 
		  __vcs_4F_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][15] .QN", 4, 
		  __vcs_50_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][6] .QN", 4, 
		  __vcs_51_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][6] .QN", 4, 
		  __vcs_52_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][13] .SI", 4, 
		  __vcs_53_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][14] .SI", 4, 
		  __vcs_54_SI_DT6vKb, "dut.DU.\\pc_current_reg[14] .SI", 3, 
		  __vcs_55_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][15] .SI", 4, 
		  __vcs_56_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][14] .QN", 4, 
		  __vcs_57_QN_DT6vKb, "dut.DU.\\pc_current_reg[15] .QN", 3, 
		  __vcs_58_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][15] .QN", 4, 
		  __vcs_59_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][13] .SI", 4, 
		  __vcs_5A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][6] .SI", 4, 
		  __vcs_5B_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][6] .SI", 4, 
		  __vcs_5C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][14] .SI", 4, 
		  __vcs_5D_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][6] .SI", 4, 
		  __vcs_5E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][6] .SI", 4, 
		  __vcs_5F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][6] .SI", 4, 
		  __vcs_60_SI_DT6vKb, "dut.DU.\\pc_current_reg[7] .SI", 3, 
		  __vcs_61_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][6] .SI", 4, 
		  __vcs_62_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][15] .SI", 4, 
		  __vcs_63_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][6] .SI", 4, 
		  __vcs_64_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][14] .QN", 4, 
		  __vcs_65_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][6] .SI", 4, 
		  __vcs_66_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][7] .QN", 4, 
		  __vcs_67_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][15] .QN", 4, 
		  __vcs_68_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][7] .QN", 4, 
		  __vcs_69_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][7] .QN", 4, 
		  __vcs_6A_QN_DT6vKb, "dut.DU.\\pc_current_reg[8] .QN", 3, 
		  __vcs_6B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][7] .QN", 4, 
		  __vcs_6C_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][7] .QN", 4, 
		  __vcs_6D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][7] .QN", 4, 
		  __vcs_6E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][7] .QN", 4, 
		  __vcs_6F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][14] .SI", 4, 
		  __vcs_70_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][15] .SI", 4, 
		  __vcs_71_SI_DT6vKb, "dut.DU.\\pc_current_reg[15] .SI", 3, 
		  __vcs_72_D_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_0/q_reg .D", 3, 
		  __vcs_73_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][15] .QN", 4, 
		  __vcs_74_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][14] .SI", 4, 
		  __vcs_75_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][7] .SI", 4, 
		  __vcs_76_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][15] .SI", 4, 
		  __vcs_77_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][7] .SI", 4, 
		  __vcs_78_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][7] .SI", 4, 
		  __vcs_79_Q_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_0/q_reg .Q", 3, 
		  __vcs_7A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][7] .SI", 4, 
		  __vcs_7B_SI_DT6vKb, "dut.DU.\\pc_current_reg[8] .SI", 3, 
		  __vcs_7C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][7] .SI", 4, 
		  __vcs_7D_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][7] .SI", 4, 
		  __vcs_7E_D_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_1/q_reg .D", 3, 
		  __vcs_7F_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][15] .QN", 4, 
		  __vcs_80_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][7] .SI", 4, 
		  __vcs_81_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][7] .SI", 4, 
		  __vcs_82_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][8] .QN", 4, 
		  __vcs_83_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][8] .QN", 4, 
		  __vcs_84_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][8] .QN", 4, 
		  __vcs_85_QN_DT6vKb, "dut.DU.\\pc_current_reg[9] .QN", 3, 
		  __vcs_86_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][8] .QN", 4, 
		  __vcs_87_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][8] .QN", 4, 
		  __vcs_88_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][8] .QN", 4, 
		  __vcs_89_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][8] .QN", 4, 
		  __vcs_8A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][15] .SI", 4, 
		  __vcs_8B_Q_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_1/q_reg .Q", 3, 
		  __vcs_8C_D_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_2/q_reg .D", 3, 
		  __vcs_8D_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][4] .Q",
		  4, __vcs_8E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][15] .SI", 4, 
		  __vcs_8F_Q_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_2/q_reg .Q", 3, 
		  __vcs_90_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][11] .Q", 4, 
		  __vcs_91_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][8] .SI", 4, 
		  __vcs_92_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][8] .Q",
		  4, __vcs_93_D_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_3/q_reg .D", 3, 
		  __vcs_94_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][8] .SI", 4, 
		  __vcs_95_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][8] .SI", 4, 
		  __vcs_96_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][8] .SI", 4, 
		  __vcs_97_SI_DT6vKb, "dut.DU.\\pc_current_reg[9] .SI", 3, 
		  __vcs_98_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][8] .SI", 4, 
		  __vcs_99_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][8] .SI", 4, 
		  __vcs_9A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][8] .SI", 4, 
		  __vcs_9B_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][8] .SI", 4, 
		  __vcs_9C_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][15] .Q", 4, 
		  __vcs_9D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][9] .QN", 4, 
		  __vcs_9E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][9] .QN", 4, 
		  __vcs_9F_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][9] .QN", 4, 
		  __vcs_A0_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][9] .QN", 4, 
		  __vcs_A1_Q_DT6vKb, 
		  "dut.snps_clk_chain_0.\\U_shftreg_0/ff_3/q_reg .Q", 3, 
		  __vcs_A2_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][9] .QN", 4, 
		  __vcs_A3_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][9] .QN", 4, 
		  __vcs_A4_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][9] .QN", 4, 
		  __vcs_A5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][10] .QN", 4, 
		  __vcs_A6_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][10] .QN", 4, 
		  __vcs_A7_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][9] .SI", 4, 
		  __vcs_A8_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][9] .SI", 4, 
		  __vcs_A9_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][9] .SI", 4, 
		  __vcs_AA_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][9] .SI", 4, 
		  __vcs_AB_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][9] .SI", 4, 
		  __vcs_AC_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][9] .SI", 4, 
		  __vcs_AD_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][9] .SI", 4, 
		  __vcs_AE_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][9] .SI", 4, 
		  __vcs_AF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][10] .SI", 4, 
		  __vcs_B0_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][10] .QN", 4, 
		  __vcs_B1_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][0] .QN", 4, 
		  __vcs_B2_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][0] .QN", 4, 
		  __vcs_B3_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][0] .QN", 4, 
		  __vcs_B4_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][0] .QN", 4, 
		  __vcs_B5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][0] .QN", 4, 
		  __vcs_B6_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][0] .QN", 4, 
		  __vcs_B7_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][0] .QN", 4, 
		  __vcs_B8_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][0] .QN", 4, 
		  __vcs_B9_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][10] .SI", 4, 
		  __vcs_BA_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][10] .QN", 4, 
		  __vcs_BB_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][11] .QN", 4, 
		  __vcs_BC_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][10] .SI", 4, 
		  __vcs_BD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][0] .SI", 4, 
		  __vcs_BE_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][0] .SI", 4, 
		  __vcs_BF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][11] .SI", 4, 
		  __vcs_C0_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][0] .SI", 4, 
		  __vcs_C1_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][10] .QN", 4, 
		  __vcs_C2_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][0] .SI", 4, 
		  __vcs_C3_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][0] .SI", 4, 
		  __vcs_C4_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][0] .SI", 4, 
		  __vcs_C5_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][0] .SI", 4, 
		  __vcs_C6_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][11] .QN", 4, 
		  __vcs_C7_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][0] .SI", 4, 
		  __vcs_C8_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][1] .QN", 4, 
		  __vcs_C9_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][12] .QN", 4, 
		  __vcs_CA_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][1] .QN", 4, 
		  __vcs_CB_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][1] .QN", 4, 
		  __vcs_CC_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][1] .QN", 4, 
		  __vcs_CD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][10] .SI", 4, 
		  __vcs_CE_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][1] .QN", 4, 
		  __vcs_CF_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][1] .QN", 4, 
		  __vcs_D0_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][1] .QN", 4, 
		  __vcs_D1_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][11] .SI", 4, 
		  __vcs_D2_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][10] .QN", 4, 
		  __vcs_D3_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][11] .QN", 4, 
		  __vcs_D4_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][12] .QN", 4, 
		  __vcs_D5_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][10] .SI", 4, 
		  __vcs_D6_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][11] .SI", 4, 
		  __vcs_D7_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][10] .QN", 4, 
		  __vcs_D8_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][1] .SI", 4, 
		  __vcs_D9_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][1] .SI", 4, 
		  __vcs_DA_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][3] .Q",
		  4, __vcs_DB_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][12] .SI", 4,
		  __vcs_DC_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][1] .SI", 4, 
		  __vcs_DD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][1] .SI", 4, 
		  __vcs_DE_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][11] .QN", 4, 
		  __vcs_DF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][1] .SI", 4, 
		  __vcs_E0_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][1] .SI", 4, 
		  __vcs_E1_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][1] .SI", 4, 
		  __vcs_E2_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][12] .QN", 4, 
		  __vcs_E3_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][1] .SI", 4, 
		  __vcs_E4_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][10] .Q", 4, 
		  __vcs_E5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][2] .QN", 4, 
		  __vcs_E6_Q_DT6vKb, "dut.DU.reg_file.\\reg_array_reg[0][7] .Q",
		  4, __vcs_E7_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][10] .SI", 4,
		  __vcs_E8_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][2] .QN", 4, 
		  __vcs_E9_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][13] .QN", 4, 
		  __vcs_EA_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][2] .QN", 4, 
		  __vcs_EB_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][2] .QN", 4, 
		  __vcs_EC_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][2] .QN", 4, 
		  __vcs_ED_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][11] .SI", 4, 
		  __vcs_EE_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][2] .QN", 4, 
		  __vcs_EF_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][10] .QN", 4, 
		  __vcs_F0_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][2] .QN", 4, 
		  __vcs_F1_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][2] .QN", 4, 
		  __vcs_F2_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][12] .SI", 4, 
		  __vcs_F3_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][14] .Q", 4, 
		  __vcs_F4_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][11] .QN", 4, 
		  __vcs_F5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][12] .QN", 4, 
		  __vcs_F6_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][10] .SI", 4, 
		  __vcs_F7_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][13] .QN", 4, 
		  __vcs_F8_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][11] .SI", 4, 
		  __vcs_F9_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][12] .SI", 4, 
		  __vcs_FA_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][11] .QN", 4, 
		  __vcs_FB_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][2] .SI", 4, 
		  __vcs_FC_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][2] .SI", 4, 
		  __vcs_FD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][2] .SI", 4, 
		  __vcs_FE_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][13] .SI", 4, 
		  __vcs_FF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][2] .SI", 4, 
		  __vcs_100_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][12] .QN", 4, 
		  __vcs_101_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][2] .SI", 4, 
		  __vcs_102_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][2] .SI", 4, 
		  __vcs_103_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][2] .SI", 4, 
		  __vcs_104_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][10] .SI", 4, 
		  __vcs_105_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][2] .SI", 4, 
		  __vcs_106_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][13] .QN", 4, 
		  __vcs_107_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][3] .QN", 4, 
		  __vcs_108_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][11] .SI", 4, 
		  __vcs_109_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][3] .QN", 4, 
		  __vcs_10A_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][14] .QN", 4, 
		  __vcs_10B_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][3] .QN", 4, 
		  __vcs_10C_QN_DT6vKb, "dut.DU.\\pc_current_reg[0] .QN", 3, 
		  __vcs_10D_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][3] .QN", 4, 
		  __vcs_10E_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][3] .QN", 4, 
		  __vcs_10F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][12] .SI", 4, 
		  __vcs_110_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][3] .QN", 4, 
		  __vcs_111_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][11] .QN", 4, 
		  __vcs_112_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][3] .QN", 4, 
		  __vcs_113_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][3] .QN", 4, 
		  __vcs_114_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][13] .SI", 4, 
		  __vcs_115_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][12] .QN", 4, 
		  __vcs_116_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][13] .QN", 4, 
		  __vcs_117_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][11] .SI", 4, 
		  __vcs_118_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][14] .QN", 4, 
		  __vcs_119_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][12] .SI", 4, 
		  __vcs_11A_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][13] .SI", 4, 
		  __vcs_11B_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][12] .QN", 4, 
		  __vcs_11C_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][3] .SI", 4, 
		  __vcs_11D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][3] .SI", 4, 
		  __vcs_11E_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][14] .SI", 4, 
		  __vcs_11F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][3] .SI", 4, 
		  __vcs_120_SI_DT6vKb, "dut.DU.\\pc_current_reg[0] .SI", 3, 
		  __vcs_121_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][13] .QN", 4, 
		  __vcs_122_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][3] .SI", 4, 
		  __vcs_123_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][3] .SI", 4, 
		  __vcs_124_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][3] .SI", 4, 
		  __vcs_125_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][11] .SI", 4, 
		  __vcs_126_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][3] .SI", 4, 
		  __vcs_127_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][0] .QN", 4, 
		  __vcs_128_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][14] .QN", 4, 
		  __vcs_129_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][3] .SI", 4, 
		  __vcs_12A_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][0] .QN", 4, 
		  __vcs_12B_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][4] .QN", 4, 
		  __vcs_12C_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][0] .QN", 4, 
		  __vcs_12D_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][4] .QN", 4, 
		  __vcs_12E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][0] .QN", 4, 
		  __vcs_12F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][12] .SI", 4, 
		  __vcs_130_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][4] .QN", 4, 
		  __vcs_131_QN_DT6vKb, "dut.DU.\\pc_current_reg[1] .QN", 3, 
		  __vcs_132_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][0] .QN", 4, 
		  __vcs_133_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][15] .QN", 4, 
		  __vcs_134_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][4] .QN", 4, 
		  __vcs_135_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][0] .QN", 4, 
		  __vcs_136_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][4] .QN", 4, 
		  __vcs_137_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][0] .QN", 4, 
		  __vcs_138_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][13] .SI", 4, 
		  __vcs_139_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][4] .QN", 4, 
		  __vcs_13A_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][0] .QN", 4, 
		  __vcs_13B_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][4] .QN", 4, 
		  __vcs_13C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][12] .QN", 4, 
		  __vcs_13D_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][4] .QN", 4, 
		  __vcs_13E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][10] .QN", 4, 
		  __vcs_13F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][14] .SI", 4, 
		  __vcs_140_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][13] .QN", 4, 
		  __vcs_141_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][14] .QN", 4, 
		  __vcs_142_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][12] .SI", 4, 
		  __vcs_143_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][15] .QN", 4, 
		  __vcs_144_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][10] .SI", 4, 
		  __vcs_145_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][13] .SI", 4, 
		  __vcs_146_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][10] .QN", 4, 
		  __vcs_147_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][0] .SI", 4, 
		  __vcs_148_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][14] .SI", 4, 
		  __vcs_149_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][13] .QN", 4, 
		  __vcs_14A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][0] .SI", 4, 
		  __vcs_14B_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][4] .SI", 4, 
		  __vcs_14C_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][0] .SI", 4, 
		  __vcs_14D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][4] .SI", 4, 
		  __vcs_14E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][0] .SI", 4, 
		  __vcs_14F_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][15] .SI", 4, 
		  __vcs_150_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][4] .SI", 4, 
		  __vcs_151_SI_DT6vKb, "dut.DU.\\pc_current_reg[1] .SI", 3, 
		  __vcs_152_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][0] .SI", 4, 
		  __vcs_153_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][4] .SI", 4, 
		  __vcs_154_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][0] .SI", 4, 
		  __vcs_155_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][14] .QN", 4, 
		  __vcs_156_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][4] .SI", 4, 
		  __vcs_157_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][0] .SI", 4, 
		  __vcs_158_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][4] .SI", 4, 
		  __vcs_159_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][0] .SI", 4, 
		  __vcs_15A_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][4] .SI", 4, 
		  __vcs_15B_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][12] .SI", 4, 
		  __vcs_15C_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][1] .QN", 4, 
		  __vcs_15D_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][15] .QN", 4, 
		  __vcs_15E_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][4] .SI", 4, 
		  __vcs_15F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][10] .SI", 4, 
		  __vcs_160_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][1] .QN", 4, 
		  __vcs_161_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][1] .QN", 4, 
		  __vcs_162_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][1] .QN", 4, 
		  __vcs_163_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][13] .SI", 4, 
		  __vcs_164_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][5] .QN", 4, 
		  __vcs_165_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][1] .QN", 4, 
		  __vcs_166_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][5] .QN", 4, 
		  __vcs_167_QN_DT6vKb, "dut.DU.\\pc_current_reg[2] .QN", 3, 
		  __vcs_168_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][1] .QN", 4, 
		  __vcs_169_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][5] .QN", 4, 
		  __vcs_16A_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][10] .QN", 4, 
		  __vcs_16B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][1] .QN", 4, 
		  __vcs_16C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][5] .QN", 4, 
		  __vcs_16D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][1] .QN", 4, 
		  __vcs_16E_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][14] .SI", 4, 
		  __vcs_16F_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][5] .QN", 4, 
		  __vcs_170_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][13] .QN", 4, 
		  __vcs_171_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][5] .QN", 4, 
		  __vcs_172_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][11] .QN", 4, 
		  __vcs_173_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][5] .QN", 4, 
		  __vcs_174_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][15] .SI", 4, 
		  __vcs_175_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][14] .QN", 4, 
		  __vcs_176_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][15] .QN", 4, 
		  __vcs_177_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][10] .SI", 4, 
		  __vcs_178_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][13] .SI", 4, 
		  __vcs_179_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][6] .Q", 4, 
		  __vcs_17A_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][11] .SI", 4, 
		  __vcs_17B_QN_DT6vKb, "dut.DU.\\pc_current_reg[10] .QN", 3, 
		  __vcs_17C_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][10] .QN", 4, 
		  __vcs_17D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][14] .SI", 4, 
		  __vcs_17E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][11] .QN", 4, 
		  __vcs_17F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][1] .SI", 4, 
		  __vcs_180_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][15] .SI", 4, 
		  __vcs_181_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][1] .SI", 4, 
		  __vcs_182_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][14] .QN", 4, 
		  __vcs_183_Q_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][13] .Q", 4, 
		  __vcs_184_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][1] .SI", 4, 
		  __vcs_185_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][5] .SI", 4, 
		  __vcs_186_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][1] .SI", 4, 
		  __vcs_187_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][5] .SI", 4, 
		  __vcs_188_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][1] .SI", 4, 
		  __vcs_189_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][5] .SI", 4, 
		  __vcs_18A_SI_DT6vKb, "dut.DU.\\pc_current_reg[2] .SI", 3, 
		  __vcs_18B_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][1] .SI", 4, 
		  __vcs_18C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][15] .QN", 4, 
		  __vcs_18D_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][5] .SI", 4, 
		  __vcs_18E_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][10] .SI", 4, 
		  __vcs_18F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][1] .SI", 4, 
		  __vcs_190_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][5] .SI", 4, 
		  __vcs_191_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][1] .SI", 4, 
		  __vcs_192_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][5] .SI", 4, 
		  __vcs_193_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][13] .SI", 4, 
		  __vcs_194_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][5] .SI", 4, 
		  __vcs_195_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][11] .SI", 4, 
		  __vcs_196_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][2] .QN", 4, 
		  __vcs_197_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][5] .SI", 4, 
		  __vcs_198_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][10] .QN", 4, 
		  __vcs_199_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][2] .QN", 4, 
		  __vcs_19A_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][6] .QN", 4, 
		  __vcs_19B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][2] .QN", 4, 
		  __vcs_19C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][6] .QN", 4, 
		  __vcs_19D_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][2] .QN", 4, 
		  __vcs_19E_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][14] .SI", 4, 
		  __vcs_19F_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][6] .QN", 4, 
		  __vcs_1A0_QN_DT6vKb, "dut.DU.\\pc_current_reg[3] .QN", 3, 
		  __vcs_1A1_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][2] .QN", 4, 
		  __vcs_1A2_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][6] .QN", 4, 
		  __vcs_1A3_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][11] .QN", 4, 
		  __vcs_1A4_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][2] .QN", 4, 
		  __vcs_1A5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][6] .QN", 4, 
		  __vcs_1A6_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][2] .QN", 4, 
		  __vcs_1A7_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][15] .SI", 4, 
		  __vcs_1A8_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][6] .QN", 4, 
		  __vcs_1A9_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][2] .QN", 4, 
		  __vcs_1AA_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][6] .QN", 4, 
		  __vcs_1AB_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][14] .QN", 4, 
		  __vcs_1AC_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][6] .QN", 4, 
		  __vcs_1AD_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][12] .QN", 4, 
		  __vcs_1AE_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][10] .SI", 4, 
		  __vcs_1AF_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][15] .QN", 4, 
		  __vcs_1B0_SI_DT6vKb, "dut.DU.\\pc_current_reg[10] .SI", 3, 
		  __vcs_1B1_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][11] .SI", 4, 
		  __vcs_1B2_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][10] .QN", 4, 
		  __vcs_1B3_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][14] .SI", 4, 
		  __vcs_1B4_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][12] .SI", 4, 
		  __vcs_1B5_QN_DT6vKb, "dut.DU.\\pc_current_reg[11] .QN", 3, 
		  __vcs_1B6_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][11] .QN", 4, 
		  __vcs_1B7_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][15] .SI", 4, 
		  __vcs_1B8_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][12] .QN", 4, 
		  __vcs_1B9_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][2] .SI", 4, 
		  __vcs_1BA_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][10] .SI", 4, 
		  __vcs_1BB_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][15] .QN", 4, 
		  __vcs_1BC_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][2] .SI", 4, 
		  __vcs_1BD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][6] .SI", 4, 
		  __vcs_1BE_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][2] .SI", 4, 
		  __vcs_1BF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][6] .SI", 4, 
		  __vcs_1C0_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][2] .SI", 4, 
		  __vcs_1C1_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][6] .SI", 4, 
		  __vcs_1C2_SI_DT6vKb, "dut.DU.\\pc_current_reg[3] .SI", 3, 
		  __vcs_1C3_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][2] .SI", 4, 
		  __vcs_1C4_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][6] .SI", 4, 
		  __vcs_1C5_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][11] .SI", 4, 
		  __vcs_1C6_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][2] .SI", 4, 
		  __vcs_1C7_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][10] .QN", 4, 
		  __vcs_1C8_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][6] .SI", 4, 
		  __vcs_1C9_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][2] .SI", 4, 
		  __vcs_1CA_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][6] .SI", 4, 
		  __vcs_1CB_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][2] .SI", 4, 
		  __vcs_1CC_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][6] .SI", 4, 
		  __vcs_1CD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][14] .SI", 4, 
		  __vcs_1CE_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][12] .SI", 4, 
		  __vcs_1CF_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][6] .SI", 4, 
		  __vcs_1D0_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][3] .QN", 4, 
		  __vcs_1D1_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][11] .QN", 4, 
		  __vcs_1D2_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][3] .QN", 4, 
		  __vcs_1D3_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][7] .QN", 4, 
		  __vcs_1D4_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][3] .QN", 4, 
		  __vcs_1D5_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][15] .SI", 4, 
		  __vcs_1D6_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][7] .QN", 4, 
		  __vcs_1D7_QN_DT6vKb, "dut.DU.\\pc_current_reg[4] .QN", 3, 
		  __vcs_1D8_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][3] .QN", 4, 
		  __vcs_1D9_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][7] .QN", 4, 
		  __vcs_1DA_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][12] .QN", 4, 
		  __vcs_1DB_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][3] .QN", 4, 
		  __vcs_1DC_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][7] .QN", 4, 
		  __vcs_1DD_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][3] .QN", 4, 
		  __vcs_1DE_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][7] .QN", 4, 
		  __vcs_1DF_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][3] .QN", 4, 
		  __vcs_1E0_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][7] .QN", 4, 
		  __vcs_1E1_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][10] .SI", 4, 
		  __vcs_1E2_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][15] .QN", 4, 
		  __vcs_1E3_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][7] .QN", 4, 
		  __vcs_1E4_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][13] .QN", 4, 
		  __vcs_1E5_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][7] .QN", 4, 
		  __vcs_1E6_SI_DT6vKb, "dut.DU.\\pc_current_reg[11] .SI", 3, 
		  __vcs_1E7_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][11] .SI", 4, 
		  __vcs_1E8_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][12] .SI", 4, 
		  __vcs_1E9_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][11] .QN", 4, 
		  __vcs_1EA_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][15] .SI", 4, 
		  __vcs_1EB_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][13] .SI", 4, 
		  __vcs_1EC_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][12] .QN", 4, 
		  __vcs_1ED_QN_DT6vKb, "dut.DU.\\pc_current_reg[12] .QN", 3, 
		  __vcs_1EE_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][10] .SI", 4, 
		  __vcs_1EF_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][13] .QN", 4, 
		  __vcs_1F0_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][3] .SI", 4, 
		  __vcs_1F1_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][3] .SI", 4, 
		  __vcs_1F2_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][11] .SI", 4, 
		  __vcs_1F3_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][3] .SI", 4, 
		  __vcs_1F4_SI_DT6vKb, "dut.DU.dm.\\memory_reg[0][7] .SI", 4, 
		  __vcs_1F5_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][3] .SI", 4, 
		  __vcs_1F6_SI_DT6vKb, "dut.DU.dm.\\memory_reg[1][7] .SI", 4, 
		  __vcs_1F7_SI_DT6vKb, "dut.DU.\\pc_current_reg[4] .SI", 3, 
		  __vcs_1F8_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][3] .SI", 4, 
		  __vcs_1F9_SI_DT6vKb, "dut.DU.dm.\\memory_reg[2][7] .SI", 4, 
		  __vcs_1FA_SI_DT6vKb, "dut.DU.dm.\\memory_reg[3][7] .SI", 4, 
		  __vcs_1FB_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][12] .SI", 4, 
		  __vcs_1FC_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][3] .SI", 4, 
		  __vcs_1FD_SI_DT6vKb, "dut.DU.dm.\\memory_reg[4][7] .SI", 4, 
		  __vcs_1FE_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][11] .QN", 4, 
		  __vcs_1FF_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][3] .SI", 4, 
		  __vcs_200_SI_DT6vKb, "dut.DU.dm.\\memory_reg[5][7] .SI", 4, 
		  __vcs_201_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][3] .SI", 4, 
		  __vcs_202_SI_DT6vKb, "dut.DU.dm.\\memory_reg[6][7] .SI", 4, 
		  __vcs_203_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][15] .SI", 4, 
		  __vcs_204_SI_DT6vKb, "dut.DU.dm.\\memory_reg[7][7] .SI", 4, 
		  __vcs_205_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][13] .SI", 4, 
		  __vcs_206_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][12] .QN", 4, 
		  __vcs_207_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][4] .QN", 4, 
		  __vcs_208_QN_DT6vKb, "dut.DU.dm.\\memory_reg[0][8] .QN", 4, 
		  __vcs_209_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][4] .QN", 4, 
		  __vcs_20A_QN_DT6vKb, "dut.DU.dm.\\memory_reg[1][8] .QN", 4, 
		  __vcs_20B_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][4] .QN", 4, 
		  __vcs_20C_QN_DT6vKb, "dut.DU.dm.\\memory_reg[2][8] .QN", 4, 
		  __vcs_20D_QN_DT6vKb, "dut.DU.\\pc_current_reg[5] .QN", 3, 
		  __vcs_20E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][4] .QN", 4, 
		  __vcs_20F_QN_DT6vKb, "dut.DU.dm.\\memory_reg[3][8] .QN", 4, 
		  __vcs_210_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[3][13] .QN", 4, 
		  __vcs_211_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][4] .QN", 4, 
		  __vcs_212_Q_DT6vKb, "dut.DU.dm.\\memory_reg[0][5] .Q", 4, 
		  __vcs_213_QN_DT6vKb, "dut.DU.dm.\\memory_reg[4][8] .QN", 4, 
		  __vcs_214_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][4] .QN", 4, 
		  __vcs_215_QN_DT6vKb, "dut.DU.dm.\\memory_reg[5][8] .QN", 4, 
		  __vcs_216_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][4] .QN", 4, 
		  __vcs_217_QN_DT6vKb, "dut.DU.dm.\\memory_reg[6][8] .QN", 4, 
		  __vcs_218_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][11] .SI", 4, 
		  __vcs_219_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][14] .QN", 4, 
		  __vcs_21A_QN_DT6vKb, "dut.DU.dm.\\memory_reg[7][8] .QN", 4, 
		  __vcs_21B_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][12] .SI", 4, 
		  __vcs_21C_SI_DT6vKb, "dut.DU.\\pc_current_reg[12] .SI", 3, 
		  __vcs_21D_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][13] .SI", 4, 
		  __vcs_21E_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[6][12] .QN", 4, 
		  __vcs_21F_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][14] .SI", 4, 
		  __vcs_220_QN_DT6vKb, "dut.DU.\\pc_current_reg[13] .QN", 3, 
		  __vcs_221_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[4][13] .QN", 4, 
		  __vcs_222_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[7][11] .SI", 4, 
		  __vcs_223_QN_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[2][14] .QN", 4, 
		  __vcs_224_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[0][4] .SI", 4, 
		  __vcs_225_Q_DT6vKb, "dut.DU.dm.\\memory_reg[0][11] .Q", 4, 
		  __vcs_226_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[1][4] .SI", 4, 
		  __vcs_227_SI_DT6vKb, 
		  "dut.DU.reg_file.\\reg_array_reg[5][12] .SI", 4);
	  $$compile_pkg(0, "", "_vcs_unit__17393910");
	end
	initial begin : DebugProcess
	  $$xmr_debugUsedPliTf("$countdrivers", "$dumpports", "$dumpportsall", 
		  "$dumpportsflush", "$dumpportslimit", "$dumpportsoff", 
		  "$dumpportson", "$fs_inject_evcd_vectors", 
		  "$fsdbAddRuntimeSignal", "$fsdbAutoSwitchDumpfile", 
		  "$fsdbDisplay", "$fsdbLog", "$fsdbSubstituteHier", 
		  "$fsdbSuppress", "$fsdbSuppressClassMethod", 
		  "$fsdbSuppressClassProp", "$fsdbSwitchDumpfile", 
		  "$fsdbTrans_add_attribute", "$fsdbTrans_add_attribute_expand",
		  "$fsdbTrans_add_relation", "$fsdbTrans_add_scope_attribute", 
		  "$fsdbTrans_add_stream_attribute", "$fsdbTrans_add_tag", 
		  "$fsdbTrans_begin", "$fsdbTrans_create_stream_begin", 
		  "$fsdbTrans_create_stream_end", "$fsdbTrans_define_attribute",
		  "$fsdbTrans_end", "$fsdbTrans_get_error_code", 
		  "$fsdbTrans_set_label", "$fsim_register_strobe", 
		  "$fsim_register_verify", "$lsi_dumpports", "$ridbDump", 
		  "$simlearn", "$sps_add_attribute", "$sps_add_relation", 
		  "$sps_begin_transaction", "$sps_create_transaction_stream", 
		  "$sps_end_transaction", "$sps_flush_file", 
		  "$sps_free_transaction", "$sps_interactive", "$sps_test", 
		  "$sps_update_label", "$vcs_get_object_id", 
		  "$vcs_get_object_type", "$vcsmemprof");
	end
endmodule

`delay_mode_path
`portcoerce
`inline
/* Source file "Risc_16_bit_netlist_scan.v", line 2844 */
`timescale 1 ns / 1 ps

(* PARTCOMP_MOD_SUFFIX = "g2J7Bb", PARTCOMP_MOD_ORIG_NAME = "Risc_16_bit" *) 

`timescale 1ns/1ps
module Risc_16_bit(clk, TEST_SI1, TEST_SI2, TEST_SI3, TEST_SI4, TEST_SE
	, TEST_SO1, TEST_SO2, TEST_SO3, TEST_SO4, scan_clk, SCAN_MODE
	, pll_bypass_2, pll_reset, test_si5, test_so5, test_si6, test_so6
	, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, test_si10
	, test_so10, test_si11, test_so11, test_si12, test_so12, test_si13
	, test_so13, test_si14, test_so14, test_si15, test_so15, test_si16
	, test_so16, test_si17, test_so17, test_si18, test_so18, test_si19
	, test_so19, test_si20, test_so20, test_si21, test_so21, test_si22
	, test_so22, test_si23, test_so23, test_si24, test_so24, test_si25
	, test_so25, test_si26, test_so26, test_si27, test_so27, test_si28
	, test_so28, test_si29, test_so29, test_si30, test_so30, test_si31
	, test_so31, test_si32, test_so32, test_si33, test_so33, test_si34
	, test_so34, test_si35, test_so35, test_si36, test_so36, test_si37
	, test_so37, test_si38, test_so38, test_si39, test_so39, test_si40
	, test_so40, test_si41, test_so41, test_si42, test_so42, test_si43
	, test_so43, test_si44, test_so44, test_si45, test_so45, test_si46
	, test_so46, test_si47, test_so47);

	input			clk;
	input			TEST_SI1;
	input			TEST_SI2;
	input			TEST_SI3;
	input			TEST_SI4;
	input			TEST_SE;
	input			scan_clk;
	input			SCAN_MODE;
	input			pll_bypass_2;
	input			pll_reset;
	input			test_si5;
	input			test_si6;
	input			test_si7;
	input			test_si8;
	input			test_si9;
	input			test_si10;
	input			test_si11;
	input			test_si12;
	input			test_si13;
	input			test_si14;
	input			test_si15;
	input			test_si16;
	input			test_si17;
	input			test_si18;
	input			test_si19;
	input			test_si20;
	input			test_si21;
	input			test_si22;
	input			test_si23;
	input			test_si24;
	input			test_si25;
	input			test_si26;
	input			test_si27;
	input			test_si28;
	input			test_si29;
	input			test_si30;
	input			test_si31;
	input			test_si32;
	input			test_si33;
	input			test_si34;
	input			test_si35;
	input			test_si36;
	input			test_si37;
	input			test_si38;
	input			test_si39;
	input			test_si40;
	input			test_si41;
	input			test_si42;
	input			test_si43;
	input			test_si44;
	input			test_si45;
	input			test_si46;
	input			test_si47;
	output			TEST_SO1;
	output			TEST_SO2;
	output			TEST_SO3;
	output			TEST_SO4;
	output			test_so5;
	output			test_so6;
	output			test_so7;
	output			test_so8;
	output			test_so9;
	output			test_so10;
	output			test_so11;
	output			test_so12;
	output			test_so13;
	output			test_so14;
	output			test_so15;
	output			test_so16;
	output			test_so17;
	output			test_so18;
	output			test_so19;
	output			test_so20;
	output			test_so21;
	output			test_so22;
	output			test_so23;
	output			test_so24;
	output			test_so25;
	output			test_so26;
	output			test_so27;
	output			test_so28;
	output			test_so29;
	output			test_so30;
	output			test_so31;
	output			test_so32;
	output			test_so33;
	output			test_so34;
	output			test_so35;
	output			test_so36;
	output			test_so37;
	output			test_so38;
	output			test_so39;
	output			test_so40;
	output			test_so41;
	output			test_so42;
	output			test_so43;
	output			test_so44;
	output			test_so45;
	output			test_so46;
	output			test_so47;
endmodule
