// Verilog netlist written by  TetraMAX(R)  U-2022.12-SP7-i20231010_191200 
// Date: Mon May 20 15:27:38 2024

module LSDNENX1 (ENB, D, Q);
input ENB, D;
output Q;
   or or0 (Q, ENB, D);
endmodule

module SDFFSSRX2 (CLK, D, RSTB, SETB, SI, SE, Q, QN);
input CLK, D, RSTB, SETB, SI, SE;
output Q, QN;
wire S, DS, D1, D2, Q_buf, setb, rstb, nD, nCLK, nSE, nSI, CLK_D_RSTB_SI_SE, RSTB_CLK_D, 
       CLK_nD_RSTB_nSI_nSE, RSTB_nCLK_D, RSTB_nCLK_nD, CLK_D_SETB_SI_SE, 
       CLK_nD_SETB_nSI_nSE, nCLK_D_SETB, nCLK_nD_SETB, D_RSTB_SI_SE, nD_RSTB_nSI_nSE, 
       CLK_D_RSTB, RSTB_CLK_nD, nCLK_D_RSTB, nCLK_nD_RSTB, D_SETB, nD_SETB, CLK_D_SETB, 
       CLK_nD_SETB, CLK_D, CLK_RSTB, CLK_SETB, CLK_nD, nCLK_D, nCLK_nD, D_SE, D_SI, D_RSTB
       , RSTB_SETB, RSTB_D_SETB, RSTB_nD_SETB, RSTB_nD, RSTB_i, SETB_i, CLK_check, D_check
       ;
reg notifier;
   pullup pullup0 (setb);
   pullup pullup1 (rstb);
   not not2 (S, SETB);
   or or3 (DS, S, D);
   and and4 (D1, DS, RSTB);
   saed90_mux saed90_mux5 (D2, D1, SI, SE);
   saed90_dff_pos saed90_dff_pos6 (Q_buf, D2, CLK, rstb, setb, notifier);
   buf buf7 (Q, Q_buf);
   not not8 (QN, Q_buf);
   not not9 (nD, D);
   not not10 (nCLK, CLK);
   not not11 (nSE, SE);
   not not12 (nSI, SI);
   and and13 (CLK_D_RSTB_SI_SE, CLK, D, RSTB, SI, SE);
   and and14 (RSTB_CLK_D, RSTB, CLK, D);
   and and15 (CLK_nD_RSTB_nSI_nSE, CLK, nD, RSTB, nSI, nSE);
   and and16 (RSTB_nCLK_D, RSTB, nCLK, D);
   and and17 (RSTB_nCLK_nD, RSTB, nCLK, nD);
   and and18 (CLK_D_SETB_SI_SE, CLK, D, SETB, SI, SE);
   and and19 (CLK_nD_SETB_nSI_nSE, CLK, nD, SETB, nSI, nSE);
   and and20 (nCLK_D_SETB, nCLK, D, SETB);
   and and21 (nCLK_nD_SETB, nCLK, nD, SETB);
   and and22 (D_RSTB_SI_SE, D, RSTB, SI, SE);
   and and23 (nD_RSTB_nSI_nSE, nD, RSTB, nSI, nSE);
   and and24 (CLK_D_RSTB, CLK, D, RSTB);
   and and25 (RSTB_CLK_nD, RSTB, CLK, nD);
   and and26 (nCLK_D_RSTB, nCLK, D, RSTB);
   and and27 (nCLK_nD_RSTB, nCLK, nD, RSTB);
   and and28 (D_SETB, D, SETB);
   and and29 (nD_SETB, nD, SETB);
   and and30 (CLK_D_SETB, CLK, D, SETB);
   and and31 (CLK_nD_SETB, CLK, nD, SETB);
   and and32 (nCLK_D_SETB, nCLK, D, SETB);
   and and33 (nCLK_nD_SETB, nCLK, nD, SETB);
   and and34 (CLK_D, CLK, D);
   and and35 (CLK_RSTB, CLK, RSTB);
   and and36 (CLK_SETB, CLK, SETB);
   and and37 (CLK_nD, CLK, nD);
   and and38 (nCLK_D, nCLK, D);
   and and39 (nCLK_nD, nCLK, nD);
   and and40 (D_SE, D, SE);
   and and41 (D_SI, D, SI);
   and and42 (D_RSTB, D, RSTB);
   and and43 (D_SETB, D, SETB);
   and and44 (RSTB_SETB, RSTB, SETB);
   and and45 (RSTB_D_SETB, RSTB, D, SETB);
   and and46 (RSTB_nD_SETB, RSTB, nD, SETB);
   and and47 (RSTB_nD, RSTB, nD);
   buf buf48 (RSTB_i, RSTB);
   buf buf49 (SETB_i, SETB);
   and and50 (CLK_check, RSTB_i, SETB_i);
   and and51 (D_check, RSTB_i, SETB_i);
endmodule

`suppress_faults
`enable_portfaults
module TIEL (ZN);
output ZN;
   buf buf0 (ZN, 1'b0);
endmodule
`disable_portfaults
`nosuppress_faults

module Instruction_Memory (pc, instruction);
input [15:0] pc;
output [15:0] instruction;
   assign instruction[0] = 1'b0;
   assign instruction[1] = 1'b0;
   assign instruction[2] = 1'b0;
   assign instruction[3] = 1'b0;
   assign instruction[4] = 1'b0;
   assign instruction[5] = 1'b0;
   assign instruction[6] = 1'b0;
   assign instruction[7] = 1'b0;
   assign instruction[8] = 1'b0;
   assign instruction[9] = 1'b0;
   assign instruction[10] = 1'b0;
   assign instruction[11] = 1'b0;
   assign instruction[12] = 1'b0;
   assign instruction[13] = 1'b0;
   assign instruction[14] = 1'b0;
   assign instruction[15] = 1'b0;
endmodule

module GPRs_test_1 (clk, reg_write_en, reg_write_dest, reg_write_data, reg_read_addr_1, 
       reg_read_data_1, reg_read_addr_2, reg_read_data_2, test_si2, test_si1, test_so2, 
       test_so1, test_se);
input clk, reg_write_en, test_si2, test_si1, test_se;
input [2:0] reg_write_dest;
input [15:0] reg_write_data;
input [2:0] reg_read_addr_1;
input [2:0] reg_read_addr_2;
output test_so2, test_so1;
output [15:0] reg_read_data_1;
output [15:0] reg_read_data_2;
wire N10, N11, N12, N13, N14, N15, \reg_array[7][15] , \reg_array[7][14] , 
       \reg_array[7][13] , \reg_array[7][12] , \reg_array[7][11] , \reg_array[7][10] , 
       \reg_array[7][9] , \reg_array[7][8] , \reg_array[7][7] , \reg_array[7][6] , 
       \reg_array[7][5] , \reg_array[7][4] , \reg_array[7][3] , \reg_array[7][2] , 
       \reg_array[7][1] , \reg_array[7][0] , \reg_array[6][15] , \reg_array[6][14] , 
       \reg_array[6][13] , \reg_array[6][12] , \reg_array[6][11] , \reg_array[6][10] , 
       \reg_array[6][9] , \reg_array[6][8] , \reg_array[6][7] , \reg_array[6][6] , 
       \reg_array[6][5] , \reg_array[6][4] , \reg_array[6][3] , \reg_array[6][2] , 
       \reg_array[6][1] , \reg_array[6][0] , \reg_array[5][15] , \reg_array[5][14] , 
       \reg_array[5][13] , \reg_array[5][12] , \reg_array[5][11] , \reg_array[5][10] , 
       \reg_array[5][9] , \reg_array[5][8] , \reg_array[5][7] , \reg_array[5][6] , 
       \reg_array[5][5] , \reg_array[5][4] , \reg_array[5][3] , \reg_array[5][2] , 
       \reg_array[5][1] , \reg_array[5][0] , \reg_array[4][15] , \reg_array[4][14] , 
       \reg_array[4][13] , \reg_array[4][12] , \reg_array[4][11] , \reg_array[4][10] , 
       \reg_array[4][9] , \reg_array[4][8] , \reg_array[4][7] , \reg_array[4][6] , 
       \reg_array[4][5] , \reg_array[4][4] , \reg_array[4][3] , \reg_array[4][2] , 
       \reg_array[4][1] , \reg_array[4][0] , \reg_array[3][15] , \reg_array[3][14] , 
       \reg_array[3][13] , \reg_array[3][12] , \reg_array[3][11] , \reg_array[3][10] , 
       \reg_array[3][9] , \reg_array[3][8] , \reg_array[3][7] , \reg_array[3][6] , 
       \reg_array[3][5] , \reg_array[3][4] , \reg_array[3][3] , \reg_array[3][2] , 
       \reg_array[3][1] , \reg_array[3][0] , \reg_array[2][15] , \reg_array[2][14] , 
       \reg_array[2][13] , \reg_array[2][12] , \reg_array[2][11] , \reg_array[2][10] , 
       \reg_array[2][9] , \reg_array[2][8] , \reg_array[2][7] , \reg_array[2][6] , 
       \reg_array[2][5] , \reg_array[2][4] , \reg_array[2][3] , \reg_array[2][2] , 
       \reg_array[2][1] , \reg_array[2][0] , \reg_array[1][15] , \reg_array[1][14] , 
       \reg_array[1][13] , \reg_array[1][12] , \reg_array[1][11] , \reg_array[1][10] , 
       \reg_array[1][9] , \reg_array[1][8] , \reg_array[1][7] , \reg_array[1][6] , 
       \reg_array[1][5] , \reg_array[1][4] , \reg_array[1][3] , \reg_array[1][2] , 
       \reg_array[1][1] , \reg_array[1][0] , \reg_array[0][15] , \reg_array[0][14] , 
       \reg_array[0][13] , \reg_array[0][12] , \reg_array[0][11] , \reg_array[0][10] , 
       \reg_array[0][9] , \reg_array[0][8] , \reg_array[0][7] , \reg_array[0][6] , 
       \reg_array[0][5] , \reg_array[0][4] , \reg_array[0][3] , \reg_array[0][2] , 
       \reg_array[0][1] , \reg_array[0][0] , n140, n141, n142, n143, n144, n145, n146, 
       n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160
       , n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
       n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187
       , n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
       n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214
       , n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
       n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241
       , n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
       n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268
       , n269, n270, n271, n272, n273, n274, n275, n276, n277, n129, n130, n131, n132, 
       n133, n134, n135, n136, n137, n138, n139, n278, n279, n280, n281, n282, n283, n284
       , n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
       n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311
       , n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
       n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338
       , n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
       n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365
       , n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
       n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392
       , n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
       n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419
       , n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
       n433, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447
       , n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
       n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474
       , n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
       n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501
       , n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
       n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528
       , n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, 
       n542, n543, n544, n545, n546, n547;
   assign N10 = reg_read_addr_1[0];
   assign N11 = reg_read_addr_1[1];
   assign N12 = reg_read_addr_1[2];
   assign N13 = reg_read_addr_2[0];
   assign N14 = reg_read_addr_2[1];
   assign N15 = reg_read_addr_2[2];
   assign test_so2 = \reg_array[7][15] ;
   assign test_so1 = \reg_array[2][5] ;
   SDFFX1 \reg_array_reg[7][15]  (.D(n277), .SI(n435), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][15] ));
   SDFFX1 \reg_array_reg[7][14]  (.D(n276), .SI(n436), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][14] ), .QN(n435));
   SDFFX1 \reg_array_reg[7][13]  (.D(n275), .SI(n437), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][13] ), .QN(n436));
   SDFFX1 \reg_array_reg[7][12]  (.D(n274), .SI(n438), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][12] ), .QN(n437));
   SDFFX1 \reg_array_reg[7][11]  (.D(n273), .SI(n439), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][11] ), .QN(n438));
   SDFFX1 \reg_array_reg[7][10]  (.D(n272), .SI(n440), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][10] ), .QN(n439));
   SDFFX1 \reg_array_reg[7][9]  (.D(n271), .SI(n441), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][9] ), .QN(n440));
   SDFFX1 \reg_array_reg[7][8]  (.D(n270), .SI(n442), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][8] ), .QN(n441));
   SDFFX1 \reg_array_reg[7][7]  (.D(n269), .SI(n443), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][7] ), .QN(n442));
   SDFFX1 \reg_array_reg[7][6]  (.D(n268), .SI(n444), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][6] ), .QN(n443));
   SDFFX1 \reg_array_reg[7][5]  (.D(n267), .SI(n445), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][5] ), .QN(n444));
   SDFFX1 \reg_array_reg[7][4]  (.D(n266), .SI(n446), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][4] ), .QN(n445));
   SDFFX1 \reg_array_reg[7][3]  (.D(n265), .SI(n447), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][3] ), .QN(n446));
   SDFFX1 \reg_array_reg[7][2]  (.D(n264), .SI(n448), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][2] ), .QN(n447));
   SDFFX1 \reg_array_reg[7][1]  (.D(n263), .SI(n449), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][1] ), .QN(n448));
   SDFFX1 \reg_array_reg[7][0]  (.D(n262), .SI(n450), .SE(test_se), .CLK(clk), .Q(
          \reg_array[7][0] ), .QN(n449));
   SDFFX1 \reg_array_reg[6][15]  (.D(n261), .SI(n451), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][15] ), .QN(n450));
   SDFFX1 \reg_array_reg[6][14]  (.D(n260), .SI(n452), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][14] ), .QN(n451));
   SDFFX1 \reg_array_reg[6][13]  (.D(n259), .SI(n453), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][13] ), .QN(n452));
   SDFFX1 \reg_array_reg[6][12]  (.D(n258), .SI(n454), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][12] ), .QN(n453));
   SDFFX1 \reg_array_reg[6][11]  (.D(n257), .SI(n455), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][11] ), .QN(n454));
   SDFFX1 \reg_array_reg[6][10]  (.D(n256), .SI(n456), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][10] ), .QN(n455));
   SDFFX1 \reg_array_reg[6][9]  (.D(n255), .SI(n457), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][9] ), .QN(n456));
   SDFFX1 \reg_array_reg[6][8]  (.D(n254), .SI(n458), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][8] ), .QN(n457));
   SDFFX1 \reg_array_reg[6][7]  (.D(n253), .SI(n459), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][7] ), .QN(n458));
   SDFFX1 \reg_array_reg[6][6]  (.D(n252), .SI(n460), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][6] ), .QN(n459));
   SDFFX1 \reg_array_reg[6][5]  (.D(n251), .SI(n461), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][5] ), .QN(n460));
   SDFFX1 \reg_array_reg[6][4]  (.D(n250), .SI(n462), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][4] ), .QN(n461));
   SDFFX1 \reg_array_reg[6][3]  (.D(n249), .SI(n463), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][3] ), .QN(n462));
   SDFFX1 \reg_array_reg[6][2]  (.D(n248), .SI(n464), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][2] ), .QN(n463));
   SDFFX1 \reg_array_reg[6][1]  (.D(n247), .SI(n465), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][1] ), .QN(n464));
   SDFFX1 \reg_array_reg[6][0]  (.D(n246), .SI(n466), .SE(test_se), .CLK(clk), .Q(
          \reg_array[6][0] ), .QN(n465));
   SDFFX1 \reg_array_reg[5][15]  (.D(n245), .SI(n467), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][15] ), .QN(n466));
   SDFFX1 \reg_array_reg[5][14]  (.D(n244), .SI(n468), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][14] ), .QN(n467));
   SDFFX1 \reg_array_reg[5][13]  (.D(n243), .SI(n469), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][13] ), .QN(n468));
   SDFFX1 \reg_array_reg[5][12]  (.D(n242), .SI(n470), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][12] ), .QN(n469));
   SDFFX1 \reg_array_reg[5][11]  (.D(n241), .SI(n471), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][11] ), .QN(n470));
   SDFFX1 \reg_array_reg[5][10]  (.D(n240), .SI(n472), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][10] ), .QN(n471));
   SDFFX1 \reg_array_reg[5][9]  (.D(n239), .SI(n473), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][9] ), .QN(n472));
   SDFFX1 \reg_array_reg[5][8]  (.D(n238), .SI(n474), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][8] ), .QN(n473));
   SDFFX1 \reg_array_reg[5][7]  (.D(n237), .SI(n475), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][7] ), .QN(n474));
   SDFFX1 \reg_array_reg[5][6]  (.D(n236), .SI(n476), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][6] ), .QN(n475));
   SDFFX1 \reg_array_reg[5][5]  (.D(n235), .SI(n477), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][5] ), .QN(n476));
   SDFFX1 \reg_array_reg[5][4]  (.D(n234), .SI(n478), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][4] ), .QN(n477));
   SDFFX1 \reg_array_reg[5][3]  (.D(n233), .SI(n479), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][3] ), .QN(n478));
   SDFFX1 \reg_array_reg[5][2]  (.D(n232), .SI(n480), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][2] ), .QN(n479));
   SDFFX1 \reg_array_reg[5][1]  (.D(n231), .SI(n481), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][1] ), .QN(n480));
   SDFFX1 \reg_array_reg[5][0]  (.D(n230), .SI(n482), .SE(test_se), .CLK(clk), .Q(
          \reg_array[5][0] ), .QN(n481));
   SDFFX1 \reg_array_reg[4][15]  (.D(n229), .SI(n483), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][15] ), .QN(n482));
   SDFFX1 \reg_array_reg[4][14]  (.D(n228), .SI(n484), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][14] ), .QN(n483));
   SDFFX1 \reg_array_reg[4][13]  (.D(n227), .SI(n485), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][13] ), .QN(n484));
   SDFFX1 \reg_array_reg[4][12]  (.D(n226), .SI(n486), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][12] ), .QN(n485));
   SDFFX1 \reg_array_reg[4][11]  (.D(n225), .SI(n487), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][11] ), .QN(n486));
   SDFFX1 \reg_array_reg[4][10]  (.D(n224), .SI(n488), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][10] ), .QN(n487));
   SDFFX1 \reg_array_reg[4][9]  (.D(n223), .SI(n489), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][9] ), .QN(n488));
   SDFFX1 \reg_array_reg[4][8]  (.D(n222), .SI(n490), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][8] ), .QN(n489));
   SDFFX1 \reg_array_reg[4][7]  (.D(n221), .SI(n491), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][7] ), .QN(n490));
   SDFFX1 \reg_array_reg[4][6]  (.D(n220), .SI(n492), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][6] ), .QN(n491));
   SDFFX1 \reg_array_reg[4][5]  (.D(n219), .SI(n493), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][5] ), .QN(n492));
   SDFFX1 \reg_array_reg[4][4]  (.D(n218), .SI(n494), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][4] ), .QN(n493));
   SDFFX1 \reg_array_reg[4][3]  (.D(n217), .SI(n495), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][3] ), .QN(n494));
   SDFFX1 \reg_array_reg[4][2]  (.D(n216), .SI(n496), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][2] ), .QN(n495));
   SDFFX1 \reg_array_reg[4][1]  (.D(n215), .SI(n497), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][1] ), .QN(n496));
   SDFFX1 \reg_array_reg[4][0]  (.D(n214), .SI(n498), .SE(test_se), .CLK(clk), .Q(
          \reg_array[4][0] ), .QN(n497));
   SDFFX1 \reg_array_reg[3][15]  (.D(n213), .SI(n499), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][15] ), .QN(n498));
   SDFFX1 \reg_array_reg[3][14]  (.D(n212), .SI(n500), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][14] ), .QN(n499));
   SDFFX1 \reg_array_reg[3][13]  (.D(n211), .SI(n501), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][13] ), .QN(n500));
   SDFFX1 \reg_array_reg[3][12]  (.D(n210), .SI(n502), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][12] ), .QN(n501));
   SDFFX1 \reg_array_reg[3][11]  (.D(n209), .SI(n503), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][11] ), .QN(n502));
   SDFFX1 \reg_array_reg[3][10]  (.D(n208), .SI(n504), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][10] ), .QN(n503));
   SDFFX1 \reg_array_reg[3][9]  (.D(n207), .SI(n505), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][9] ), .QN(n504));
   SDFFX1 \reg_array_reg[3][8]  (.D(n206), .SI(n506), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][8] ), .QN(n505));
   SDFFX1 \reg_array_reg[3][7]  (.D(n205), .SI(n507), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][7] ), .QN(n506));
   SDFFX1 \reg_array_reg[3][6]  (.D(n204), .SI(n508), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][6] ), .QN(n507));
   SDFFX1 \reg_array_reg[3][5]  (.D(n203), .SI(n509), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][5] ), .QN(n508));
   SDFFX1 \reg_array_reg[3][4]  (.D(n202), .SI(n510), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][4] ), .QN(n509));
   SDFFX1 \reg_array_reg[3][3]  (.D(n201), .SI(n511), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][3] ), .QN(n510));
   SDFFX1 \reg_array_reg[3][2]  (.D(n200), .SI(n512), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][2] ), .QN(n511));
   SDFFX1 \reg_array_reg[3][1]  (.D(n199), .SI(n513), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][1] ), .QN(n512));
   SDFFX1 \reg_array_reg[3][0]  (.D(n198), .SI(n514), .SE(test_se), .CLK(clk), .Q(
          \reg_array[3][0] ), .QN(n513));
   SDFFX1 \reg_array_reg[2][15]  (.D(n197), .SI(n515), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][15] ), .QN(n514));
   SDFFX1 \reg_array_reg[2][14]  (.D(n196), .SI(n516), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][14] ), .QN(n515));
   SDFFX1 \reg_array_reg[2][13]  (.D(n195), .SI(n517), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][13] ), .QN(n516));
   SDFFX1 \reg_array_reg[2][12]  (.D(n194), .SI(n518), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][12] ), .QN(n517));
   SDFFX1 \reg_array_reg[2][11]  (.D(n193), .SI(n519), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][11] ), .QN(n518));
   SDFFX1 \reg_array_reg[2][10]  (.D(n192), .SI(n520), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][10] ), .QN(n519));
   SDFFX1 \reg_array_reg[2][9]  (.D(n191), .SI(n521), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][9] ), .QN(n520));
   SDFFX1 \reg_array_reg[2][8]  (.D(n190), .SI(n522), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][8] ), .QN(n521));
   SDFFX1 \reg_array_reg[2][7]  (.D(n189), .SI(n523), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][7] ), .QN(n522));
   SDFFX1 \reg_array_reg[2][6]  (.D(n188), .SI(test_si2), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][6] ), .QN(n523));
   SDFFX1 \reg_array_reg[2][5]  (.D(n187), .SI(n524), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][5] ));
   SDFFX1 \reg_array_reg[2][4]  (.D(n186), .SI(n525), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][4] ), .QN(n524));
   SDFFX1 \reg_array_reg[2][3]  (.D(n185), .SI(n526), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][3] ), .QN(n525));
   SDFFX1 \reg_array_reg[2][2]  (.D(n184), .SI(n527), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][2] ), .QN(n526));
   SDFFX1 \reg_array_reg[2][1]  (.D(n183), .SI(n528), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][1] ), .QN(n527));
   SDFFX1 \reg_array_reg[2][0]  (.D(n182), .SI(n529), .SE(test_se), .CLK(clk), .Q(
          \reg_array[2][0] ), .QN(n528));
   SDFFX1 \reg_array_reg[1][15]  (.D(n181), .SI(n530), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][15] ), .QN(n529));
   SDFFX1 \reg_array_reg[1][14]  (.D(n180), .SI(n531), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][14] ), .QN(n530));
   SDFFX1 \reg_array_reg[1][13]  (.D(n179), .SI(n532), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][13] ), .QN(n531));
   SDFFX1 \reg_array_reg[1][12]  (.D(n178), .SI(n533), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][12] ), .QN(n532));
   SDFFX1 \reg_array_reg[1][11]  (.D(n177), .SI(n534), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][11] ), .QN(n533));
   SDFFX1 \reg_array_reg[1][10]  (.D(n176), .SI(n535), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][10] ), .QN(n534));
   SDFFX1 \reg_array_reg[1][9]  (.D(n175), .SI(n536), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][9] ), .QN(n535));
   SDFFX1 \reg_array_reg[1][8]  (.D(n174), .SI(n537), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][8] ), .QN(n536));
   SDFFX1 \reg_array_reg[1][7]  (.D(n173), .SI(n538), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][7] ), .QN(n537));
   SDFFX1 \reg_array_reg[1][6]  (.D(n172), .SI(n539), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][6] ), .QN(n538));
   SDFFX1 \reg_array_reg[1][5]  (.D(n171), .SI(n540), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][5] ), .QN(n539));
   SDFFX1 \reg_array_reg[1][4]  (.D(n170), .SI(n541), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][4] ), .QN(n540));
   SDFFX1 \reg_array_reg[1][3]  (.D(n169), .SI(n542), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][3] ), .QN(n541));
   SDFFX1 \reg_array_reg[1][2]  (.D(n168), .SI(n543), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][2] ), .QN(n542));
   SDFFX1 \reg_array_reg[1][1]  (.D(n167), .SI(n544), .SE(test_se), .CLK(clk), .Q(
          \reg_array[1][1] ), .QN(n543));
   SDFFX1 \reg_array_reg[1][0]  (.D(n166), .SI(\reg_array[0][15] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[1][0] ), .QN(n544));
   SDFFX1 \reg_array_reg[0][15]  (.D(n165), .SI(\reg_array[0][14] ), .SE(test_se), .CLK(
          clk), .Q(\reg_array[0][15] ));
   SDFFX1 \reg_array_reg[0][14]  (.D(n164), .SI(\reg_array[0][13] ), .SE(test_se), .CLK(
          clk), .Q(\reg_array[0][14] ));
   SDFFX1 \reg_array_reg[0][13]  (.D(n163), .SI(\reg_array[0][12] ), .SE(test_se), .CLK(
          clk), .Q(\reg_array[0][13] ));
   SDFFX1 \reg_array_reg[0][12]  (.D(n162), .SI(\reg_array[0][11] ), .SE(test_se), .CLK(
          clk), .Q(\reg_array[0][12] ));
   SDFFX1 \reg_array_reg[0][11]  (.D(n161), .SI(\reg_array[0][10] ), .SE(test_se), .CLK(
          clk), .Q(\reg_array[0][11] ));
   SDFFX1 \reg_array_reg[0][10]  (.D(n160), .SI(\reg_array[0][9] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][10] ));
   SDFFX1 \reg_array_reg[0][9]  (.D(n159), .SI(\reg_array[0][8] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][9] ));
   SDFFX1 \reg_array_reg[0][8]  (.D(n158), .SI(\reg_array[0][7] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][8] ));
   SDFFX1 \reg_array_reg[0][7]  (.D(n157), .SI(\reg_array[0][6] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][7] ));
   SDFFX1 \reg_array_reg[0][6]  (.D(n156), .SI(\reg_array[0][5] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][6] ));
   SDFFX1 \reg_array_reg[0][5]  (.D(n155), .SI(\reg_array[0][4] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][5] ));
   SDFFX1 \reg_array_reg[0][4]  (.D(n154), .SI(\reg_array[0][3] ), .SE(test_se), .CLK(clk)
          , .Q(\reg_array[0][4] ));
   SDFFX1 \reg_array_reg[0][3]  (.D(n153), .SI(n545), .SE(test_se), .CLK(clk), .Q(
          \reg_array[0][3] ));
   SDFFX1 \reg_array_reg[0][2]  (.D(n152), .SI(n546), .SE(test_se), .CLK(clk), .Q(
          \reg_array[0][2] ), .QN(n545));
   SDFFX1 \reg_array_reg[0][1]  (.D(n151), .SI(n547), .SE(test_se), .CLK(clk), .Q(
          \reg_array[0][1] ), .QN(n546));
   SDFFX1 \reg_array_reg[0][0]  (.D(n150), .SI(test_si1), .SE(test_se), .CLK(clk), .Q(
          \reg_array[0][0] ), .QN(n547));
   AO22X1 U142 (.IN1(reg_write_data[0]), .IN2(n426), .IN3(\reg_array[0][0] ), .IN4(n140), .
          Q(n150));
   AO22X1 U143 (.IN1(reg_write_data[1]), .IN2(n426), .IN3(\reg_array[0][1] ), .IN4(n140), .
          Q(n151));
   AO22X1 U144 (.IN1(reg_write_data[2]), .IN2(n426), .IN3(\reg_array[0][2] ), .IN4(n140), .
          Q(n152));
   AO22X1 U145 (.IN1(reg_write_data[3]), .IN2(n426), .IN3(\reg_array[0][3] ), .IN4(n140), .
          Q(n153));
   AO22X1 U146 (.IN1(reg_write_data[4]), .IN2(n426), .IN3(\reg_array[0][4] ), .IN4(n140), .
          Q(n154));
   AO22X1 U147 (.IN1(reg_write_data[5]), .IN2(n426), .IN3(\reg_array[0][5] ), .IN4(n140), .
          Q(n155));
   AO22X1 U148 (.IN1(reg_write_data[6]), .IN2(n426), .IN3(\reg_array[0][6] ), .IN4(n140), .
          Q(n156));
   AO22X1 U149 (.IN1(reg_write_data[7]), .IN2(n426), .IN3(\reg_array[0][7] ), .IN4(n140), .
          Q(n157));
   AO22X1 U150 (.IN1(reg_write_data[8]), .IN2(n426), .IN3(\reg_array[0][8] ), .IN4(n140), .
          Q(n158));
   AO22X1 U151 (.IN1(reg_write_data[9]), .IN2(n426), .IN3(\reg_array[0][9] ), .IN4(n140), .
          Q(n159));
   AO22X1 U152 (.IN1(reg_write_data[10]), .IN2(n426), .IN3(\reg_array[0][10] ), .IN4(n140)
          , .Q(n160));
   AO22X1 U153 (.IN1(reg_write_data[11]), .IN2(n426), .IN3(\reg_array[0][11] ), .IN4(n140)
          , .Q(n161));
   AO22X1 U154 (.IN1(reg_write_data[12]), .IN2(n426), .IN3(\reg_array[0][12] ), .IN4(n140)
          , .Q(n162));
   AO22X1 U155 (.IN1(reg_write_data[13]), .IN2(n426), .IN3(\reg_array[0][13] ), .IN4(n140)
          , .Q(n163));
   AO22X1 U156 (.IN1(reg_write_data[14]), .IN2(n426), .IN3(\reg_array[0][14] ), .IN4(n140)
          , .Q(n164));
   AO22X1 U157 (.IN1(reg_write_data[15]), .IN2(n426), .IN3(\reg_array[0][15] ), .IN4(n140)
          , .Q(n165));
   AO22X1 U159 (.IN1(n428), .IN2(reg_write_data[0]), .IN3(\reg_array[1][0] ), .IN4(n142), .
          Q(n166));
   AO22X1 U160 (.IN1(n428), .IN2(reg_write_data[1]), .IN3(\reg_array[1][1] ), .IN4(n142), .
          Q(n167));
   AO22X1 U161 (.IN1(n428), .IN2(reg_write_data[2]), .IN3(\reg_array[1][2] ), .IN4(n142), .
          Q(n168));
   AO22X1 U162 (.IN1(n428), .IN2(reg_write_data[3]), .IN3(\reg_array[1][3] ), .IN4(n142), .
          Q(n169));
   AO22X1 U163 (.IN1(n428), .IN2(reg_write_data[4]), .IN3(\reg_array[1][4] ), .IN4(n142), .
          Q(n170));
   AO22X1 U164 (.IN1(n428), .IN2(reg_write_data[5]), .IN3(\reg_array[1][5] ), .IN4(n142), .
          Q(n171));
   AO22X1 U165 (.IN1(n428), .IN2(reg_write_data[6]), .IN3(\reg_array[1][6] ), .IN4(n142), .
          Q(n172));
   AO22X1 U166 (.IN1(n428), .IN2(reg_write_data[7]), .IN3(\reg_array[1][7] ), .IN4(n142), .
          Q(n173));
   AO22X1 U167 (.IN1(n428), .IN2(reg_write_data[8]), .IN3(\reg_array[1][8] ), .IN4(n142), .
          Q(n174));
   AO22X1 U168 (.IN1(n428), .IN2(reg_write_data[9]), .IN3(\reg_array[1][9] ), .IN4(n142), .
          Q(n175));
   AO22X1 U169 (.IN1(n428), .IN2(reg_write_data[10]), .IN3(\reg_array[1][10] ), .IN4(n142)
          , .Q(n176));
   AO22X1 U170 (.IN1(n428), .IN2(reg_write_data[11]), .IN3(\reg_array[1][11] ), .IN4(n142)
          , .Q(n177));
   AO22X1 U171 (.IN1(n428), .IN2(reg_write_data[12]), .IN3(\reg_array[1][12] ), .IN4(n142)
          , .Q(n178));
   AO22X1 U172 (.IN1(n428), .IN2(reg_write_data[13]), .IN3(\reg_array[1][13] ), .IN4(n142)
          , .Q(n179));
   AO22X1 U173 (.IN1(n428), .IN2(reg_write_data[14]), .IN3(\reg_array[1][14] ), .IN4(n142)
          , .Q(n180));
   AO22X1 U174 (.IN1(n428), .IN2(reg_write_data[15]), .IN3(\reg_array[1][15] ), .IN4(n142)
          , .Q(n181));
   AO22X1 U176 (.IN1(n425), .IN2(reg_write_data[0]), .IN3(\reg_array[2][0] ), .IN4(n143), .
          Q(n182));
   AO22X1 U177 (.IN1(n425), .IN2(reg_write_data[1]), .IN3(\reg_array[2][1] ), .IN4(n143), .
          Q(n183));
   AO22X1 U178 (.IN1(n425), .IN2(reg_write_data[2]), .IN3(\reg_array[2][2] ), .IN4(n143), .
          Q(n184));
   AO22X1 U179 (.IN1(n425), .IN2(reg_write_data[3]), .IN3(\reg_array[2][3] ), .IN4(n143), .
          Q(n185));
   AO22X1 U180 (.IN1(n425), .IN2(reg_write_data[4]), .IN3(\reg_array[2][4] ), .IN4(n143), .
          Q(n186));
   AO22X1 U181 (.IN1(n425), .IN2(reg_write_data[5]), .IN3(\reg_array[2][5] ), .IN4(n143), .
          Q(n187));
   AO22X1 U182 (.IN1(n425), .IN2(reg_write_data[6]), .IN3(\reg_array[2][6] ), .IN4(n143), .
          Q(n188));
   AO22X1 U183 (.IN1(n425), .IN2(reg_write_data[7]), .IN3(\reg_array[2][7] ), .IN4(n143), .
          Q(n189));
   AO22X1 U184 (.IN1(n425), .IN2(reg_write_data[8]), .IN3(\reg_array[2][8] ), .IN4(n143), .
          Q(n190));
   AO22X1 U185 (.IN1(n425), .IN2(reg_write_data[9]), .IN3(\reg_array[2][9] ), .IN4(n143), .
          Q(n191));
   AO22X1 U186 (.IN1(n425), .IN2(reg_write_data[10]), .IN3(\reg_array[2][10] ), .IN4(n143)
          , .Q(n192));
   AO22X1 U187 (.IN1(n425), .IN2(reg_write_data[11]), .IN3(\reg_array[2][11] ), .IN4(n143)
          , .Q(n193));
   AO22X1 U188 (.IN1(n425), .IN2(reg_write_data[12]), .IN3(\reg_array[2][12] ), .IN4(n143)
          , .Q(n194));
   AO22X1 U189 (.IN1(n425), .IN2(reg_write_data[13]), .IN3(\reg_array[2][13] ), .IN4(n143)
          , .Q(n195));
   AO22X1 U190 (.IN1(n425), .IN2(reg_write_data[14]), .IN3(\reg_array[2][14] ), .IN4(n143)
          , .Q(n196));
   AO22X1 U191 (.IN1(n425), .IN2(reg_write_data[15]), .IN3(\reg_array[2][15] ), .IN4(n143)
          , .Q(n197));
   AO22X1 U193 (.IN1(n429), .IN2(reg_write_data[0]), .IN3(\reg_array[3][0] ), .IN4(n144), .
          Q(n198));
   AO22X1 U194 (.IN1(n429), .IN2(reg_write_data[1]), .IN3(\reg_array[3][1] ), .IN4(n144), .
          Q(n199));
   AO22X1 U195 (.IN1(n429), .IN2(reg_write_data[2]), .IN3(\reg_array[3][2] ), .IN4(n144), .
          Q(n200));
   AO22X1 U196 (.IN1(n429), .IN2(reg_write_data[3]), .IN3(\reg_array[3][3] ), .IN4(n144), .
          Q(n201));
   AO22X1 U197 (.IN1(n429), .IN2(reg_write_data[4]), .IN3(\reg_array[3][4] ), .IN4(n144), .
          Q(n202));
   AO22X1 U198 (.IN1(n429), .IN2(reg_write_data[5]), .IN3(\reg_array[3][5] ), .IN4(n144), .
          Q(n203));
   AO22X1 U199 (.IN1(n429), .IN2(reg_write_data[6]), .IN3(\reg_array[3][6] ), .IN4(n144), .
          Q(n204));
   AO22X1 U200 (.IN1(n429), .IN2(reg_write_data[7]), .IN3(\reg_array[3][7] ), .IN4(n144), .
          Q(n205));
   AO22X1 U201 (.IN1(n429), .IN2(reg_write_data[8]), .IN3(\reg_array[3][8] ), .IN4(n144), .
          Q(n206));
   AO22X1 U202 (.IN1(n429), .IN2(reg_write_data[9]), .IN3(\reg_array[3][9] ), .IN4(n144), .
          Q(n207));
   AO22X1 U203 (.IN1(n429), .IN2(reg_write_data[10]), .IN3(\reg_array[3][10] ), .IN4(n144)
          , .Q(n208));
   AO22X1 U204 (.IN1(n429), .IN2(reg_write_data[11]), .IN3(\reg_array[3][11] ), .IN4(n144)
          , .Q(n209));
   AO22X1 U205 (.IN1(n429), .IN2(reg_write_data[12]), .IN3(\reg_array[3][12] ), .IN4(n144)
          , .Q(n210));
   AO22X1 U206 (.IN1(n429), .IN2(reg_write_data[13]), .IN3(\reg_array[3][13] ), .IN4(n144)
          , .Q(n211));
   AO22X1 U207 (.IN1(n429), .IN2(reg_write_data[14]), .IN3(\reg_array[3][14] ), .IN4(n144)
          , .Q(n212));
   AO22X1 U208 (.IN1(n429), .IN2(reg_write_data[15]), .IN3(\reg_array[3][15] ), .IN4(n144)
          , .Q(n213));
   AO22X1 U210 (.IN1(n424), .IN2(reg_write_data[0]), .IN3(\reg_array[4][0] ), .IN4(n145), .
          Q(n214));
   AO22X1 U211 (.IN1(n424), .IN2(reg_write_data[1]), .IN3(\reg_array[4][1] ), .IN4(n145), .
          Q(n215));
   AO22X1 U212 (.IN1(n424), .IN2(reg_write_data[2]), .IN3(\reg_array[4][2] ), .IN4(n145), .
          Q(n216));
   AO22X1 U213 (.IN1(n424), .IN2(reg_write_data[3]), .IN3(\reg_array[4][3] ), .IN4(n145), .
          Q(n217));
   AO22X1 U214 (.IN1(n424), .IN2(reg_write_data[4]), .IN3(\reg_array[4][4] ), .IN4(n145), .
          Q(n218));
   AO22X1 U215 (.IN1(n424), .IN2(reg_write_data[5]), .IN3(\reg_array[4][5] ), .IN4(n145), .
          Q(n219));
   AO22X1 U216 (.IN1(n424), .IN2(reg_write_data[6]), .IN3(\reg_array[4][6] ), .IN4(n145), .
          Q(n220));
   AO22X1 U217 (.IN1(n424), .IN2(reg_write_data[7]), .IN3(\reg_array[4][7] ), .IN4(n145), .
          Q(n221));
   AO22X1 U218 (.IN1(n424), .IN2(reg_write_data[8]), .IN3(\reg_array[4][8] ), .IN4(n145), .
          Q(n222));
   AO22X1 U219 (.IN1(n424), .IN2(reg_write_data[9]), .IN3(\reg_array[4][9] ), .IN4(n145), .
          Q(n223));
   AO22X1 U220 (.IN1(n424), .IN2(reg_write_data[10]), .IN3(\reg_array[4][10] ), .IN4(n145)
          , .Q(n224));
   AO22X1 U221 (.IN1(n424), .IN2(reg_write_data[11]), .IN3(\reg_array[4][11] ), .IN4(n145)
          , .Q(n225));
   AO22X1 U222 (.IN1(n424), .IN2(reg_write_data[12]), .IN3(\reg_array[4][12] ), .IN4(n145)
          , .Q(n226));
   AO22X1 U223 (.IN1(n424), .IN2(reg_write_data[13]), .IN3(\reg_array[4][13] ), .IN4(n145)
          , .Q(n227));
   AO22X1 U224 (.IN1(n424), .IN2(reg_write_data[14]), .IN3(\reg_array[4][14] ), .IN4(n145)
          , .Q(n228));
   AO22X1 U225 (.IN1(n424), .IN2(reg_write_data[15]), .IN3(\reg_array[4][15] ), .IN4(n145)
          , .Q(n229));
   AO22X1 U227 (.IN1(n430), .IN2(reg_write_data[0]), .IN3(\reg_array[5][0] ), .IN4(n147), .
          Q(n230));
   AO22X1 U228 (.IN1(n430), .IN2(reg_write_data[1]), .IN3(\reg_array[5][1] ), .IN4(n147), .
          Q(n231));
   AO22X1 U229 (.IN1(n430), .IN2(reg_write_data[2]), .IN3(\reg_array[5][2] ), .IN4(n147), .
          Q(n232));
   AO22X1 U230 (.IN1(n430), .IN2(reg_write_data[3]), .IN3(\reg_array[5][3] ), .IN4(n147), .
          Q(n233));
   AO22X1 U231 (.IN1(n430), .IN2(reg_write_data[4]), .IN3(\reg_array[5][4] ), .IN4(n147), .
          Q(n234));
   AO22X1 U232 (.IN1(n430), .IN2(reg_write_data[5]), .IN3(\reg_array[5][5] ), .IN4(n147), .
          Q(n235));
   AO22X1 U233 (.IN1(n430), .IN2(reg_write_data[6]), .IN3(\reg_array[5][6] ), .IN4(n147), .
          Q(n236));
   AO22X1 U234 (.IN1(n430), .IN2(reg_write_data[7]), .IN3(\reg_array[5][7] ), .IN4(n147), .
          Q(n237));
   AO22X1 U235 (.IN1(n430), .IN2(reg_write_data[8]), .IN3(\reg_array[5][8] ), .IN4(n147), .
          Q(n238));
   AO22X1 U236 (.IN1(n430), .IN2(reg_write_data[9]), .IN3(\reg_array[5][9] ), .IN4(n147), .
          Q(n239));
   AO22X1 U237 (.IN1(n430), .IN2(reg_write_data[10]), .IN3(\reg_array[5][10] ), .IN4(n147)
          , .Q(n240));
   AO22X1 U238 (.IN1(n430), .IN2(reg_write_data[11]), .IN3(\reg_array[5][11] ), .IN4(n147)
          , .Q(n241));
   AO22X1 U239 (.IN1(n430), .IN2(reg_write_data[12]), .IN3(\reg_array[5][12] ), .IN4(n147)
          , .Q(n242));
   AO22X1 U240 (.IN1(n430), .IN2(reg_write_data[13]), .IN3(\reg_array[5][13] ), .IN4(n147)
          , .Q(n243));
   AO22X1 U241 (.IN1(n430), .IN2(reg_write_data[14]), .IN3(\reg_array[5][14] ), .IN4(n147)
          , .Q(n244));
   AO22X1 U242 (.IN1(n430), .IN2(reg_write_data[15]), .IN3(\reg_array[5][15] ), .IN4(n147)
          , .Q(n245));
   AO22X1 U244 (.IN1(n423), .IN2(reg_write_data[0]), .IN3(\reg_array[6][0] ), .IN4(n148), .
          Q(n246));
   AO22X1 U245 (.IN1(n423), .IN2(reg_write_data[1]), .IN3(\reg_array[6][1] ), .IN4(n148), .
          Q(n247));
   AO22X1 U246 (.IN1(n423), .IN2(reg_write_data[2]), .IN3(\reg_array[6][2] ), .IN4(n148), .
          Q(n248));
   AO22X1 U247 (.IN1(n423), .IN2(reg_write_data[3]), .IN3(\reg_array[6][3] ), .IN4(n148), .
          Q(n249));
   AO22X1 U248 (.IN1(n423), .IN2(reg_write_data[4]), .IN3(\reg_array[6][4] ), .IN4(n148), .
          Q(n250));
   AO22X1 U249 (.IN1(n423), .IN2(reg_write_data[5]), .IN3(\reg_array[6][5] ), .IN4(n148), .
          Q(n251));
   AO22X1 U250 (.IN1(n423), .IN2(reg_write_data[6]), .IN3(\reg_array[6][6] ), .IN4(n148), .
          Q(n252));
   AO22X1 U251 (.IN1(n423), .IN2(reg_write_data[7]), .IN3(\reg_array[6][7] ), .IN4(n148), .
          Q(n253));
   AO22X1 U252 (.IN1(n423), .IN2(reg_write_data[8]), .IN3(\reg_array[6][8] ), .IN4(n148), .
          Q(n254));
   AO22X1 U253 (.IN1(n423), .IN2(reg_write_data[9]), .IN3(\reg_array[6][9] ), .IN4(n148), .
          Q(n255));
   AO22X1 U254 (.IN1(n423), .IN2(reg_write_data[10]), .IN3(\reg_array[6][10] ), .IN4(n148)
          , .Q(n256));
   AO22X1 U255 (.IN1(n423), .IN2(reg_write_data[11]), .IN3(\reg_array[6][11] ), .IN4(n148)
          , .Q(n257));
   AO22X1 U256 (.IN1(n423), .IN2(reg_write_data[12]), .IN3(\reg_array[6][12] ), .IN4(n148)
          , .Q(n258));
   AO22X1 U257 (.IN1(n423), .IN2(reg_write_data[13]), .IN3(\reg_array[6][13] ), .IN4(n148)
          , .Q(n259));
   AO22X1 U258 (.IN1(n423), .IN2(reg_write_data[14]), .IN3(\reg_array[6][14] ), .IN4(n148)
          , .Q(n260));
   AO22X1 U259 (.IN1(n423), .IN2(reg_write_data[15]), .IN3(\reg_array[6][15] ), .IN4(n148)
          , .Q(n261));
   AO22X1 U261 (.IN1(n431), .IN2(reg_write_data[0]), .IN3(\reg_array[7][0] ), .IN4(n149), .
          Q(n262));
   AO22X1 U262 (.IN1(n431), .IN2(reg_write_data[1]), .IN3(\reg_array[7][1] ), .IN4(n149), .
          Q(n263));
   AO22X1 U263 (.IN1(n431), .IN2(reg_write_data[2]), .IN3(\reg_array[7][2] ), .IN4(n149), .
          Q(n264));
   AO22X1 U264 (.IN1(n431), .IN2(reg_write_data[3]), .IN3(\reg_array[7][3] ), .IN4(n149), .
          Q(n265));
   AO22X1 U265 (.IN1(n431), .IN2(reg_write_data[4]), .IN3(\reg_array[7][4] ), .IN4(n149), .
          Q(n266));
   AO22X1 U266 (.IN1(n431), .IN2(reg_write_data[5]), .IN3(\reg_array[7][5] ), .IN4(n149), .
          Q(n267));
   AO22X1 U267 (.IN1(n431), .IN2(reg_write_data[6]), .IN3(\reg_array[7][6] ), .IN4(n149), .
          Q(n268));
   AO22X1 U268 (.IN1(n431), .IN2(reg_write_data[7]), .IN3(\reg_array[7][7] ), .IN4(n149), .
          Q(n269));
   AO22X1 U269 (.IN1(n431), .IN2(reg_write_data[8]), .IN3(\reg_array[7][8] ), .IN4(n149), .
          Q(n270));
   AO22X1 U270 (.IN1(n431), .IN2(reg_write_data[9]), .IN3(\reg_array[7][9] ), .IN4(n149), .
          Q(n271));
   AO22X1 U271 (.IN1(n431), .IN2(reg_write_data[10]), .IN3(\reg_array[7][10] ), .IN4(n149)
          , .Q(n272));
   AO22X1 U272 (.IN1(n431), .IN2(reg_write_data[11]), .IN3(\reg_array[7][11] ), .IN4(n149)
          , .Q(n273));
   AO22X1 U273 (.IN1(n431), .IN2(reg_write_data[12]), .IN3(\reg_array[7][12] ), .IN4(n149)
          , .Q(n274));
   AO22X1 U274 (.IN1(n431), .IN2(reg_write_data[13]), .IN3(\reg_array[7][13] ), .IN4(n149)
          , .Q(n275));
   AO22X1 U275 (.IN1(n431), .IN2(reg_write_data[14]), .IN3(\reg_array[7][14] ), .IN4(n149)
          , .Q(n276));
   AO22X1 U276 (.IN1(n431), .IN2(reg_write_data[15]), .IN3(\reg_array[7][15] ), .IN4(n149)
          , .Q(n277));
   AND2X1 U278 (.IN1(reg_write_dest[2]), .IN2(reg_write_en), .Q(n146));
   INVX0 U130 (.INP(n140), .ZN(n426));
   INVX0 U131 (.INP(n145), .ZN(n424));
   INVX0 U132 (.INP(n142), .ZN(n428));
   INVX0 U133 (.INP(n143), .ZN(n425));
   INVX0 U134 (.INP(n144), .ZN(n429));
   INVX0 U135 (.INP(n147), .ZN(n430));
   INVX0 U136 (.INP(n148), .ZN(n423));
   INVX0 U137 (.INP(n149), .ZN(n431));
   AND2X1 U138 (.IN1(n131), .IN2(n344), .Q(n334));
   AND2X1 U139 (.IN1(n347), .IN2(n422), .Q(n412));
   AND2X1 U140 (.IN1(n133), .IN2(n344), .Q(n331));
   AND2X1 U141 (.IN1(n349), .IN2(n422), .Q(n409));
   NAND3X0 U158 (.IN1(n427), .IN2(n432), .IN3(n141), .QN(n140));
   NAND3X0 U175 (.IN1(n427), .IN2(n432), .IN3(n146), .QN(n145));
   AND2X1 U192 (.IN1(n130), .IN2(n344), .Q(n335));
   AND2X1 U209 (.IN1(n346), .IN2(n422), .Q(n413));
   AND2X1 U226 (.IN1(n132), .IN2(n344), .Q(n332));
   AND2X1 U243 (.IN1(n348), .IN2(n422), .Q(n410));
   AND2X1 U260 (.IN1(n131), .IN2(N10), .Q(n339));
   AND2X1 U277 (.IN1(n347), .IN2(N13), .Q(n417));
   AND2X1 U279 (.IN1(n133), .IN2(N10), .Q(n336));
   AND2X1 U280 (.IN1(n349), .IN2(N13), .Q(n414));
   NAND3X0 U281 (.IN1(reg_write_dest[0]), .IN2(n432), .IN3(n146), .QN(n147));
   NAND3X0 U282 (.IN1(reg_write_dest[1]), .IN2(n427), .IN3(n146), .QN(n148));
   NAND3X0 U283 (.IN1(reg_write_dest[1]), .IN2(reg_write_dest[0]), .IN3(n146), .QN(n149)
          );
   NAND3X0 U284 (.IN1(reg_write_dest[0]), .IN2(n141), .IN3(reg_write_dest[1]), .QN(n144)
          );
   NAND3X0 U285 (.IN1(n141), .IN2(n432), .IN3(reg_write_dest[0]), .QN(n142));
   NAND3X0 U286 (.IN1(n141), .IN2(n427), .IN3(reg_write_dest[1]), .QN(n143));
   AND2X1 U287 (.IN1(n130), .IN2(N10), .Q(n340));
   AND2X1 U288 (.IN1(n346), .IN2(N13), .Q(n418));
   AND2X1 U289 (.IN1(N10), .IN2(n132), .Q(n337));
   AND2X1 U290 (.IN1(N13), .IN2(n348), .Q(n415));
   NOR2X0 U291 (.IN1(n433), .IN2(reg_write_dest[2]), .QN(n141));
   INVX0 U292 (.INP(reg_write_en), .ZN(n433));
   INVX0 U293 (.INP(N10), .ZN(n344));
   INVX0 U294 (.INP(N13), .ZN(n422));
   INVX0 U295 (.INP(reg_write_dest[1]), .ZN(n432));
   INVX0 U296 (.INP(reg_write_dest[0]), .ZN(n427));
   INVX0 U297 (.INP(N11), .ZN(n343));
   INVX0 U298 (.INP(N14), .ZN(n421));
   NOR2X0 U299 (.IN1(N11), .IN2(N12), .QN(n130));
   NOR2X0 U300 (.IN1(n343), .IN2(N12), .QN(n131));
   AND2X1 U301 (.IN1(N12), .IN2(N11), .Q(n132));
   AND2X1 U302 (.IN1(N12), .IN2(n343), .Q(n133));
   AO22X1 U303 (.IN1(\reg_array[6][0] ), .IN2(n332), .IN3(\reg_array[4][0] ), .IN4(n331), .
          Q(n129));
   AO221X1 U304 (.IN1(\reg_array[0][0] ), .IN2(n335), .IN3(\reg_array[2][0] ), .IN4(n334)
          , .IN5(n129), .Q(n136));
   AO22X1 U305 (.IN1(\reg_array[7][0] ), .IN2(n337), .IN3(\reg_array[5][0] ), .IN4(n336), .
          Q(n134));
   AO221X1 U306 (.IN1(\reg_array[1][0] ), .IN2(n340), .IN3(\reg_array[3][0] ), .IN4(n339)
          , .IN5(n134), .Q(n135));
   OR2X1 U307 (.IN1(n136), .IN2(n135), .Q(reg_read_data_1[0]));
   AO22X1 U308 (.IN1(\reg_array[6][1] ), .IN2(n332), .IN3(\reg_array[4][1] ), .IN4(n331), .
          Q(n137));
   AO221X1 U309 (.IN1(\reg_array[0][1] ), .IN2(n335), .IN3(\reg_array[2][1] ), .IN4(n334)
          , .IN5(n137), .Q(n278));
   AO22X1 U310 (.IN1(\reg_array[7][1] ), .IN2(n337), .IN3(\reg_array[5][1] ), .IN4(n336), .
          Q(n138));
   AO221X1 U311 (.IN1(\reg_array[1][1] ), .IN2(n340), .IN3(\reg_array[3][1] ), .IN4(n339)
          , .IN5(n138), .Q(n139));
   OR2X1 U312 (.IN1(n278), .IN2(n139), .Q(reg_read_data_1[1]));
   AO22X1 U313 (.IN1(\reg_array[6][2] ), .IN2(n332), .IN3(\reg_array[4][2] ), .IN4(n331), .
          Q(n279));
   AO221X1 U314 (.IN1(\reg_array[0][2] ), .IN2(n335), .IN3(\reg_array[2][2] ), .IN4(n334)
          , .IN5(n279), .Q(n282));
   AO22X1 U315 (.IN1(\reg_array[7][2] ), .IN2(n337), .IN3(\reg_array[5][2] ), .IN4(n336), .
          Q(n280));
   AO221X1 U316 (.IN1(\reg_array[1][2] ), .IN2(n340), .IN3(\reg_array[3][2] ), .IN4(n339)
          , .IN5(n280), .Q(n281));
   OR2X1 U317 (.IN1(n282), .IN2(n281), .Q(reg_read_data_1[2]));
   AO22X1 U318 (.IN1(\reg_array[6][3] ), .IN2(n332), .IN3(\reg_array[4][3] ), .IN4(n331), .
          Q(n283));
   AO221X1 U319 (.IN1(\reg_array[0][3] ), .IN2(n335), .IN3(\reg_array[2][3] ), .IN4(n334)
          , .IN5(n283), .Q(n286));
   AO22X1 U320 (.IN1(\reg_array[7][3] ), .IN2(n337), .IN3(\reg_array[5][3] ), .IN4(n336), .
          Q(n284));
   AO221X1 U321 (.IN1(\reg_array[1][3] ), .IN2(n340), .IN3(\reg_array[3][3] ), .IN4(n339)
          , .IN5(n284), .Q(n285));
   OR2X1 U322 (.IN1(n286), .IN2(n285), .Q(reg_read_data_1[3]));
   AO22X1 U323 (.IN1(\reg_array[6][4] ), .IN2(n332), .IN3(\reg_array[4][4] ), .IN4(n331), .
          Q(n287));
   AO221X1 U324 (.IN1(\reg_array[0][4] ), .IN2(n335), .IN3(\reg_array[2][4] ), .IN4(n334)
          , .IN5(n287), .Q(n290));
   AO22X1 U325 (.IN1(\reg_array[7][4] ), .IN2(n337), .IN3(\reg_array[5][4] ), .IN4(n336), .
          Q(n288));
   AO221X1 U326 (.IN1(\reg_array[1][4] ), .IN2(n340), .IN3(\reg_array[3][4] ), .IN4(n339)
          , .IN5(n288), .Q(n289));
   OR2X1 U327 (.IN1(n290), .IN2(n289), .Q(reg_read_data_1[4]));
   AO22X1 U328 (.IN1(\reg_array[6][5] ), .IN2(n332), .IN3(\reg_array[4][5] ), .IN4(n331), .
          Q(n291));
   AO221X1 U329 (.IN1(\reg_array[0][5] ), .IN2(n335), .IN3(\reg_array[2][5] ), .IN4(n334)
          , .IN5(n291), .Q(n294));
   AO22X1 U330 (.IN1(\reg_array[7][5] ), .IN2(n337), .IN3(\reg_array[5][5] ), .IN4(n336), .
          Q(n292));
   AO221X1 U331 (.IN1(\reg_array[1][5] ), .IN2(n340), .IN3(\reg_array[3][5] ), .IN4(n339)
          , .IN5(n292), .Q(n293));
   OR2X1 U332 (.IN1(n294), .IN2(n293), .Q(reg_read_data_1[5]));
   AO22X1 U333 (.IN1(\reg_array[6][6] ), .IN2(n332), .IN3(\reg_array[4][6] ), .IN4(n331), .
          Q(n295));
   AO221X1 U334 (.IN1(\reg_array[0][6] ), .IN2(n335), .IN3(\reg_array[2][6] ), .IN4(n334)
          , .IN5(n295), .Q(n298));
   AO22X1 U335 (.IN1(\reg_array[7][6] ), .IN2(n337), .IN3(\reg_array[5][6] ), .IN4(n336), .
          Q(n296));
   AO221X1 U336 (.IN1(\reg_array[1][6] ), .IN2(n340), .IN3(\reg_array[3][6] ), .IN4(n339)
          , .IN5(n296), .Q(n297));
   OR2X1 U337 (.IN1(n298), .IN2(n297), .Q(reg_read_data_1[6]));
   AO22X1 U338 (.IN1(\reg_array[6][7] ), .IN2(n332), .IN3(\reg_array[4][7] ), .IN4(n331), .
          Q(n299));
   AO221X1 U339 (.IN1(\reg_array[0][7] ), .IN2(n335), .IN3(\reg_array[2][7] ), .IN4(n334)
          , .IN5(n299), .Q(n302));
   AO22X1 U340 (.IN1(\reg_array[7][7] ), .IN2(n337), .IN3(\reg_array[5][7] ), .IN4(n336), .
          Q(n300));
   AO221X1 U341 (.IN1(\reg_array[1][7] ), .IN2(n340), .IN3(\reg_array[3][7] ), .IN4(n339)
          , .IN5(n300), .Q(n301));
   OR2X1 U342 (.IN1(n302), .IN2(n301), .Q(reg_read_data_1[7]));
   AO22X1 U343 (.IN1(\reg_array[6][8] ), .IN2(n332), .IN3(\reg_array[4][8] ), .IN4(n331), .
          Q(n303));
   AO221X1 U344 (.IN1(\reg_array[0][8] ), .IN2(n335), .IN3(\reg_array[2][8] ), .IN4(n334)
          , .IN5(n303), .Q(n306));
   AO22X1 U345 (.IN1(\reg_array[7][8] ), .IN2(n337), .IN3(\reg_array[5][8] ), .IN4(n336), .
          Q(n304));
   AO221X1 U346 (.IN1(\reg_array[1][8] ), .IN2(n340), .IN3(\reg_array[3][8] ), .IN4(n339)
          , .IN5(n304), .Q(n305));
   OR2X1 U347 (.IN1(n306), .IN2(n305), .Q(reg_read_data_1[8]));
   AO22X1 U348 (.IN1(\reg_array[6][9] ), .IN2(n332), .IN3(\reg_array[4][9] ), .IN4(n331), .
          Q(n307));
   AO221X1 U349 (.IN1(\reg_array[0][9] ), .IN2(n335), .IN3(\reg_array[2][9] ), .IN4(n334)
          , .IN5(n307), .Q(n310));
   AO22X1 U350 (.IN1(\reg_array[7][9] ), .IN2(n337), .IN3(\reg_array[5][9] ), .IN4(n336), .
          Q(n308));
   AO221X1 U351 (.IN1(\reg_array[1][9] ), .IN2(n340), .IN3(\reg_array[3][9] ), .IN4(n339)
          , .IN5(n308), .Q(n309));
   OR2X1 U352 (.IN1(n310), .IN2(n309), .Q(reg_read_data_1[9]));
   AO22X1 U353 (.IN1(\reg_array[6][10] ), .IN2(n332), .IN3(\reg_array[4][10] ), .IN4(n331)
          , .Q(n311));
   AO221X1 U354 (.IN1(\reg_array[0][10] ), .IN2(n335), .IN3(\reg_array[2][10] ), .IN4(n334)
          , .IN5(n311), .Q(n314));
   AO22X1 U355 (.IN1(\reg_array[7][10] ), .IN2(n337), .IN3(\reg_array[5][10] ), .IN4(n336)
          , .Q(n312));
   AO221X1 U356 (.IN1(\reg_array[1][10] ), .IN2(n340), .IN3(\reg_array[3][10] ), .IN4(n339)
          , .IN5(n312), .Q(n313));
   OR2X1 U357 (.IN1(n314), .IN2(n313), .Q(reg_read_data_1[10]));
   AO22X1 U358 (.IN1(\reg_array[6][11] ), .IN2(n332), .IN3(\reg_array[4][11] ), .IN4(n331)
          , .Q(n315));
   AO221X1 U359 (.IN1(\reg_array[0][11] ), .IN2(n335), .IN3(\reg_array[2][11] ), .IN4(n334)
          , .IN5(n315), .Q(n318));
   AO22X1 U360 (.IN1(\reg_array[7][11] ), .IN2(n337), .IN3(\reg_array[5][11] ), .IN4(n336)
          , .Q(n316));
   AO221X1 U361 (.IN1(\reg_array[1][11] ), .IN2(n340), .IN3(\reg_array[3][11] ), .IN4(n339)
          , .IN5(n316), .Q(n317));
   OR2X1 U362 (.IN1(n318), .IN2(n317), .Q(reg_read_data_1[11]));
   AO22X1 U363 (.IN1(\reg_array[6][12] ), .IN2(n332), .IN3(\reg_array[4][12] ), .IN4(n331)
          , .Q(n319));
   AO221X1 U364 (.IN1(\reg_array[0][12] ), .IN2(n335), .IN3(\reg_array[2][12] ), .IN4(n334)
          , .IN5(n319), .Q(n322));
   AO22X1 U365 (.IN1(\reg_array[7][12] ), .IN2(n337), .IN3(\reg_array[5][12] ), .IN4(n336)
          , .Q(n320));
   AO221X1 U366 (.IN1(\reg_array[1][12] ), .IN2(n340), .IN3(\reg_array[3][12] ), .IN4(n339)
          , .IN5(n320), .Q(n321));
   OR2X1 U367 (.IN1(n322), .IN2(n321), .Q(reg_read_data_1[12]));
   AO22X1 U368 (.IN1(\reg_array[6][13] ), .IN2(n332), .IN3(\reg_array[4][13] ), .IN4(n331)
          , .Q(n323));
   AO221X1 U369 (.IN1(\reg_array[0][13] ), .IN2(n335), .IN3(\reg_array[2][13] ), .IN4(n334)
          , .IN5(n323), .Q(n326));
   AO22X1 U370 (.IN1(\reg_array[7][13] ), .IN2(n337), .IN3(\reg_array[5][13] ), .IN4(n336)
          , .Q(n324));
   AO221X1 U371 (.IN1(\reg_array[1][13] ), .IN2(n340), .IN3(\reg_array[3][13] ), .IN4(n339)
          , .IN5(n324), .Q(n325));
   OR2X1 U372 (.IN1(n326), .IN2(n325), .Q(reg_read_data_1[13]));
   AO22X1 U373 (.IN1(\reg_array[6][14] ), .IN2(n332), .IN3(\reg_array[4][14] ), .IN4(n331)
          , .Q(n327));
   AO221X1 U374 (.IN1(\reg_array[0][14] ), .IN2(n335), .IN3(\reg_array[2][14] ), .IN4(n334)
          , .IN5(n327), .Q(n330));
   AO22X1 U375 (.IN1(\reg_array[7][14] ), .IN2(n337), .IN3(\reg_array[5][14] ), .IN4(n336)
          , .Q(n328));
   AO221X1 U376 (.IN1(\reg_array[1][14] ), .IN2(n340), .IN3(\reg_array[3][14] ), .IN4(n339)
          , .IN5(n328), .Q(n329));
   OR2X1 U377 (.IN1(n330), .IN2(n329), .Q(reg_read_data_1[14]));
   AO22X1 U378 (.IN1(\reg_array[6][15] ), .IN2(n332), .IN3(\reg_array[4][15] ), .IN4(n331)
          , .Q(n333));
   AO221X1 U379 (.IN1(\reg_array[0][15] ), .IN2(n335), .IN3(\reg_array[2][15] ), .IN4(n334)
          , .IN5(n333), .Q(n342));
   AO22X1 U380 (.IN1(\reg_array[7][15] ), .IN2(n337), .IN3(\reg_array[5][15] ), .IN4(n336)
          , .Q(n338));
   AO221X1 U381 (.IN1(\reg_array[1][15] ), .IN2(n340), .IN3(\reg_array[3][15] ), .IN4(n339)
          , .IN5(n338), .Q(n341));
   OR2X1 U382 (.IN1(n342), .IN2(n341), .Q(reg_read_data_1[15]));
   NOR2X0 U383 (.IN1(N14), .IN2(N15), .QN(n346));
   NOR2X0 U384 (.IN1(n421), .IN2(N15), .QN(n347));
   AND2X1 U385 (.IN1(N15), .IN2(N14), .Q(n348));
   AND2X1 U386 (.IN1(N15), .IN2(n421), .Q(n349));
   AO22X1 U387 (.IN1(\reg_array[6][0] ), .IN2(n410), .IN3(\reg_array[4][0] ), .IN4(n409), .
          Q(n345));
   AO221X1 U388 (.IN1(\reg_array[0][0] ), .IN2(n413), .IN3(\reg_array[2][0] ), .IN4(n412)
          , .IN5(n345), .Q(n352));
   AO22X1 U389 (.IN1(\reg_array[7][0] ), .IN2(n415), .IN3(\reg_array[5][0] ), .IN4(n414), .
          Q(n350));
   AO221X1 U390 (.IN1(\reg_array[1][0] ), .IN2(n418), .IN3(\reg_array[3][0] ), .IN4(n417)
          , .IN5(n350), .Q(n351));
   OR2X1 U391 (.IN1(n352), .IN2(n351), .Q(reg_read_data_2[0]));
   AO22X1 U392 (.IN1(\reg_array[6][1] ), .IN2(n410), .IN3(\reg_array[4][1] ), .IN4(n409), .
          Q(n353));
   AO221X1 U393 (.IN1(\reg_array[0][1] ), .IN2(n413), .IN3(\reg_array[2][1] ), .IN4(n412)
          , .IN5(n353), .Q(n356));
   AO22X1 U394 (.IN1(\reg_array[7][1] ), .IN2(n415), .IN3(\reg_array[5][1] ), .IN4(n414), .
          Q(n354));
   AO221X1 U395 (.IN1(\reg_array[1][1] ), .IN2(n418), .IN3(\reg_array[3][1] ), .IN4(n417)
          , .IN5(n354), .Q(n355));
   OR2X1 U396 (.IN1(n356), .IN2(n355), .Q(reg_read_data_2[1]));
   AO22X1 U397 (.IN1(\reg_array[6][2] ), .IN2(n410), .IN3(\reg_array[4][2] ), .IN4(n409), .
          Q(n357));
   AO221X1 U398 (.IN1(\reg_array[0][2] ), .IN2(n413), .IN3(\reg_array[2][2] ), .IN4(n412)
          , .IN5(n357), .Q(n360));
   AO22X1 U399 (.IN1(\reg_array[7][2] ), .IN2(n415), .IN3(\reg_array[5][2] ), .IN4(n414), .
          Q(n358));
   AO221X1 U400 (.IN1(\reg_array[1][2] ), .IN2(n418), .IN3(\reg_array[3][2] ), .IN4(n417)
          , .IN5(n358), .Q(n359));
   OR2X1 U401 (.IN1(n360), .IN2(n359), .Q(reg_read_data_2[2]));
   AO22X1 U402 (.IN1(\reg_array[6][3] ), .IN2(n410), .IN3(\reg_array[4][3] ), .IN4(n409), .
          Q(n361));
   AO221X1 U403 (.IN1(\reg_array[0][3] ), .IN2(n413), .IN3(\reg_array[2][3] ), .IN4(n412)
          , .IN5(n361), .Q(n364));
   AO22X1 U404 (.IN1(\reg_array[7][3] ), .IN2(n415), .IN3(\reg_array[5][3] ), .IN4(n414), .
          Q(n362));
   AO221X1 U405 (.IN1(\reg_array[1][3] ), .IN2(n418), .IN3(\reg_array[3][3] ), .IN4(n417)
          , .IN5(n362), .Q(n363));
   OR2X1 U406 (.IN1(n364), .IN2(n363), .Q(reg_read_data_2[3]));
   AO22X1 U407 (.IN1(\reg_array[6][4] ), .IN2(n410), .IN3(\reg_array[4][4] ), .IN4(n409), .
          Q(n365));
   AO221X1 U408 (.IN1(\reg_array[0][4] ), .IN2(n413), .IN3(\reg_array[2][4] ), .IN4(n412)
          , .IN5(n365), .Q(n368));
   AO22X1 U409 (.IN1(\reg_array[7][4] ), .IN2(n415), .IN3(\reg_array[5][4] ), .IN4(n414), .
          Q(n366));
   AO221X1 U410 (.IN1(\reg_array[1][4] ), .IN2(n418), .IN3(\reg_array[3][4] ), .IN4(n417)
          , .IN5(n366), .Q(n367));
   OR2X1 U411 (.IN1(n368), .IN2(n367), .Q(reg_read_data_2[4]));
   AO22X1 U412 (.IN1(\reg_array[6][5] ), .IN2(n410), .IN3(\reg_array[4][5] ), .IN4(n409), .
          Q(n369));
   AO221X1 U413 (.IN1(\reg_array[0][5] ), .IN2(n413), .IN3(\reg_array[2][5] ), .IN4(n412)
          , .IN5(n369), .Q(n372));
   AO22X1 U414 (.IN1(\reg_array[7][5] ), .IN2(n415), .IN3(\reg_array[5][5] ), .IN4(n414), .
          Q(n370));
   AO221X1 U415 (.IN1(\reg_array[1][5] ), .IN2(n418), .IN3(\reg_array[3][5] ), .IN4(n417)
          , .IN5(n370), .Q(n371));
   OR2X1 U416 (.IN1(n372), .IN2(n371), .Q(reg_read_data_2[5]));
   AO22X1 U417 (.IN1(\reg_array[6][6] ), .IN2(n410), .IN3(\reg_array[4][6] ), .IN4(n409), .
          Q(n373));
   AO221X1 U418 (.IN1(\reg_array[0][6] ), .IN2(n413), .IN3(\reg_array[2][6] ), .IN4(n412)
          , .IN5(n373), .Q(n376));
   AO22X1 U419 (.IN1(\reg_array[7][6] ), .IN2(n415), .IN3(\reg_array[5][6] ), .IN4(n414), .
          Q(n374));
   AO221X1 U420 (.IN1(\reg_array[1][6] ), .IN2(n418), .IN3(\reg_array[3][6] ), .IN4(n417)
          , .IN5(n374), .Q(n375));
   OR2X1 U421 (.IN1(n376), .IN2(n375), .Q(reg_read_data_2[6]));
   AO22X1 U422 (.IN1(\reg_array[6][7] ), .IN2(n410), .IN3(\reg_array[4][7] ), .IN4(n409), .
          Q(n377));
   AO221X1 U423 (.IN1(\reg_array[0][7] ), .IN2(n413), .IN3(\reg_array[2][7] ), .IN4(n412)
          , .IN5(n377), .Q(n380));
   AO22X1 U424 (.IN1(\reg_array[7][7] ), .IN2(n415), .IN3(\reg_array[5][7] ), .IN4(n414), .
          Q(n378));
   AO221X1 U425 (.IN1(\reg_array[1][7] ), .IN2(n418), .IN3(\reg_array[3][7] ), .IN4(n417)
          , .IN5(n378), .Q(n379));
   OR2X1 U426 (.IN1(n380), .IN2(n379), .Q(reg_read_data_2[7]));
   AO22X1 U427 (.IN1(\reg_array[6][8] ), .IN2(n410), .IN3(\reg_array[4][8] ), .IN4(n409), .
          Q(n381));
   AO221X1 U428 (.IN1(\reg_array[0][8] ), .IN2(n413), .IN3(\reg_array[2][8] ), .IN4(n412)
          , .IN5(n381), .Q(n384));
   AO22X1 U429 (.IN1(\reg_array[7][8] ), .IN2(n415), .IN3(\reg_array[5][8] ), .IN4(n414), .
          Q(n382));
   AO221X1 U430 (.IN1(\reg_array[1][8] ), .IN2(n418), .IN3(\reg_array[3][8] ), .IN4(n417)
          , .IN5(n382), .Q(n383));
   OR2X1 U431 (.IN1(n384), .IN2(n383), .Q(reg_read_data_2[8]));
   AO22X1 U432 (.IN1(\reg_array[6][9] ), .IN2(n410), .IN3(\reg_array[4][9] ), .IN4(n409), .
          Q(n385));
   AO221X1 U433 (.IN1(\reg_array[0][9] ), .IN2(n413), .IN3(\reg_array[2][9] ), .IN4(n412)
          , .IN5(n385), .Q(n388));
   AO22X1 U434 (.IN1(\reg_array[7][9] ), .IN2(n415), .IN3(\reg_array[5][9] ), .IN4(n414), .
          Q(n386));
   AO221X1 U435 (.IN1(\reg_array[1][9] ), .IN2(n418), .IN3(\reg_array[3][9] ), .IN4(n417)
          , .IN5(n386), .Q(n387));
   OR2X1 U436 (.IN1(n388), .IN2(n387), .Q(reg_read_data_2[9]));
   AO22X1 U437 (.IN1(\reg_array[6][10] ), .IN2(n410), .IN3(\reg_array[4][10] ), .IN4(n409)
          , .Q(n389));
   AO221X1 U438 (.IN1(\reg_array[0][10] ), .IN2(n413), .IN3(\reg_array[2][10] ), .IN4(n412)
          , .IN5(n389), .Q(n392));
   AO22X1 U439 (.IN1(\reg_array[7][10] ), .IN2(n415), .IN3(\reg_array[5][10] ), .IN4(n414)
          , .Q(n390));
   AO221X1 U440 (.IN1(\reg_array[1][10] ), .IN2(n418), .IN3(\reg_array[3][10] ), .IN4(n417)
          , .IN5(n390), .Q(n391));
   OR2X1 U441 (.IN1(n392), .IN2(n391), .Q(reg_read_data_2[10]));
   AO22X1 U442 (.IN1(\reg_array[6][11] ), .IN2(n410), .IN3(\reg_array[4][11] ), .IN4(n409)
          , .Q(n393));
   AO221X1 U443 (.IN1(\reg_array[0][11] ), .IN2(n413), .IN3(\reg_array[2][11] ), .IN4(n412)
          , .IN5(n393), .Q(n396));
   AO22X1 U444 (.IN1(\reg_array[7][11] ), .IN2(n415), .IN3(\reg_array[5][11] ), .IN4(n414)
          , .Q(n394));
   AO221X1 U445 (.IN1(\reg_array[1][11] ), .IN2(n418), .IN3(\reg_array[3][11] ), .IN4(n417)
          , .IN5(n394), .Q(n395));
   OR2X1 U446 (.IN1(n396), .IN2(n395), .Q(reg_read_data_2[11]));
   AO22X1 U447 (.IN1(\reg_array[6][12] ), .IN2(n410), .IN3(\reg_array[4][12] ), .IN4(n409)
          , .Q(n397));
   AO221X1 U448 (.IN1(\reg_array[0][12] ), .IN2(n413), .IN3(\reg_array[2][12] ), .IN4(n412)
          , .IN5(n397), .Q(n400));
   AO22X1 U449 (.IN1(\reg_array[7][12] ), .IN2(n415), .IN3(\reg_array[5][12] ), .IN4(n414)
          , .Q(n398));
   AO221X1 U450 (.IN1(\reg_array[1][12] ), .IN2(n418), .IN3(\reg_array[3][12] ), .IN4(n417)
          , .IN5(n398), .Q(n399));
   OR2X1 U451 (.IN1(n400), .IN2(n399), .Q(reg_read_data_2[12]));
   AO22X1 U452 (.IN1(\reg_array[6][13] ), .IN2(n410), .IN3(\reg_array[4][13] ), .IN4(n409)
          , .Q(n401));
   AO221X1 U453 (.IN1(\reg_array[0][13] ), .IN2(n413), .IN3(\reg_array[2][13] ), .IN4(n412)
          , .IN5(n401), .Q(n404));
   AO22X1 U454 (.IN1(\reg_array[7][13] ), .IN2(n415), .IN3(\reg_array[5][13] ), .IN4(n414)
          , .Q(n402));
   AO221X1 U455 (.IN1(\reg_array[1][13] ), .IN2(n418), .IN3(\reg_array[3][13] ), .IN4(n417)
          , .IN5(n402), .Q(n403));
   OR2X1 U456 (.IN1(n404), .IN2(n403), .Q(reg_read_data_2[13]));
   AO22X1 U457 (.IN1(\reg_array[6][14] ), .IN2(n410), .IN3(\reg_array[4][14] ), .IN4(n409)
          , .Q(n405));
   AO221X1 U458 (.IN1(\reg_array[0][14] ), .IN2(n413), .IN3(\reg_array[2][14] ), .IN4(n412)
          , .IN5(n405), .Q(n408));
   AO22X1 U459 (.IN1(\reg_array[7][14] ), .IN2(n415), .IN3(\reg_array[5][14] ), .IN4(n414)
          , .Q(n406));
   AO221X1 U460 (.IN1(\reg_array[1][14] ), .IN2(n418), .IN3(\reg_array[3][14] ), .IN4(n417)
          , .IN5(n406), .Q(n407));
   OR2X1 U461 (.IN1(n408), .IN2(n407), .Q(reg_read_data_2[14]));
   AO22X1 U462 (.IN1(\reg_array[6][15] ), .IN2(n410), .IN3(\reg_array[4][15] ), .IN4(n409)
          , .Q(n411));
   AO221X1 U463 (.IN1(\reg_array[0][15] ), .IN2(n413), .IN3(\reg_array[2][15] ), .IN4(n412)
          , .IN5(n411), .Q(n420));
   AO22X1 U464 (.IN1(\reg_array[7][15] ), .IN2(n415), .IN3(\reg_array[5][15] ), .IN4(n414)
          , .Q(n416));
   AO221X1 U465 (.IN1(\reg_array[1][15] ), .IN2(n418), .IN3(\reg_array[3][15] ), .IN4(n417)
          , .IN5(n416), .Q(n419));
   OR2X1 U466 (.IN1(n420), .IN2(n419), .Q(reg_read_data_2[15]));
endmodule

module alu_control (ALU_Control, ALUOp, Function);
input [1:0] ALUOp;
input [3:0] Function;
output [2:0] ALU_Control;
wire n5, n6, n7, n8, n9, n10, n11, n12, n1, n2, n3, n4;
   NOR3X0 U10 (.IN1(n5), .IN2(n6), .IN3(n7), .QN(ALU_Control[2]));
   OA22X1 U11 (.IN1(n8), .IN2(n9), .IN3(n2), .IN4(n4), .Q(n6));
   NOR3X0 U12 (.IN1(n10), .IN2(Function[1]), .IN3(n5), .QN(ALU_Control[1]));
   OR2X1 U13 (.IN1(ALUOp[0]), .IN2(ALUOp[1]), .Q(n5));
   XOR2X1 U14 (.IN1(n4), .IN2(Function[2]), .Q(n10));
   NOR3X0 U15 (.IN1(n1), .IN2(n2), .IN3(n12), .QN(n11));
   XOR2X1 U16 (.IN1(n4), .IN2(n7), .Q(n12));
   XOR2X1 U17 (.IN1(Function[1]), .IN2(Function[2]), .Q(n7));
   NAND2X1 U3 (.IN1(n1), .IN2(n4), .QN(n9));
   OA21X1 U4 (.IN1(ALUOp[0]), .IN2(n11), .IN3(n3), .Q(ALU_Control[0]));
   INVX0 U5 (.INP(ALUOp[1]), .ZN(n3));
   INVX0 U6 (.INP(n8), .ZN(n2));
   INVX0 U7 (.INP(Function[3]), .ZN(n4));
   INVX0 U8 (.INP(Function[0]), .ZN(n1));
   NAND2X1 U9 (.IN1(Function[2]), .IN2(Function[1]), .QN(n8));
endmodule

module ALU_DW01_sub_0 (A, B, CI, DIFF, CO);
input CI;
input [15:0] A;
input [15:0] B;
output CO;
output [15:0] DIFF;
wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16;
wire [16:0] carry;
   FADDX1 U2_14 (.A(A[14]), .B(n5), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]));
   FADDX1 U2_13 (.A(A[13]), .B(n6), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]));
   FADDX1 U2_12 (.A(A[12]), .B(n7), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]));
   FADDX1 U2_11 (.A(A[11]), .B(n8), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]));
   FADDX1 U2_10 (.A(A[10]), .B(n9), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]));
   FADDX1 U2_9 (.A(A[9]), .B(n10), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]));
   FADDX1 U2_8 (.A(A[8]), .B(n11), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]));
   FADDX1 U2_7 (.A(A[7]), .B(n12), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]));
   FADDX1 U2_6 (.A(A[6]), .B(n13), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]));
   FADDX1 U2_5 (.A(A[5]), .B(n14), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]));
   FADDX1 U2_4 (.A(A[4]), .B(n3), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]));
   FADDX1 U2_3 (.A(A[3]), .B(n2), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]));
   FADDX1 U2_2 (.A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]));
   FADDX1 U2_1 (.A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]));
   XOR3X1 U2_15 (.IN1(A[15]), .IN2(n4), .IN3(carry[15]), .Q(DIFF[15]));
   INVX0 U1 (.INP(B[15]), .ZN(n4));
   INVX0 U2 (.INP(B[6]), .ZN(n13));
   INVX0 U3 (.INP(B[2]), .ZN(n15));
   INVX0 U4 (.INP(B[4]), .ZN(n3));
   INVX0 U5 (.INP(B[8]), .ZN(n11));
   INVX0 U6 (.INP(B[10]), .ZN(n9));
   INVX0 U7 (.INP(B[12]), .ZN(n7));
   INVX0 U8 (.INP(B[14]), .ZN(n5));
   NAND2X1 U9 (.IN1(n1), .IN2(B[0]), .QN(carry[1]));
   INVX0 U10 (.INP(B[1]), .ZN(n16));
   INVX0 U11 (.INP(A[0]), .ZN(n1));
   INVX0 U12 (.INP(B[3]), .ZN(n2));
   INVX0 U13 (.INP(B[7]), .ZN(n12));
   INVX0 U14 (.INP(B[9]), .ZN(n10));
   INVX0 U15 (.INP(B[11]), .ZN(n8));
   INVX0 U16 (.INP(B[5]), .ZN(n14));
   INVX0 U17 (.INP(B[13]), .ZN(n6));
   XOR2X1 U18 (.IN1(B[0]), .IN2(A[0]), .Q(DIFF[0]));
endmodule

module ALU_DW01_add_0_DW01_add_2 (A, B, CI, SUM, CO);
input CI;
input [15:0] A;
input [15:0] B;
output CO;
output [15:0] SUM;
wire n1;
wire [15:1] carry;
   FADDX1 U1_14 (.A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(SUM[14]));
   FADDX1 U1_13 (.A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(SUM[13]));
   FADDX1 U1_12 (.A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(SUM[12]));
   FADDX1 U1_11 (.A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(SUM[11]));
   FADDX1 U1_10 (.A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(SUM[10]));
   FADDX1 U1_9 (.A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]));
   FADDX1 U1_8 (.A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]));
   FADDX1 U1_7 (.A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]));
   FADDX1 U1_6 (.A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]));
   FADDX1 U1_5 (.A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]));
   FADDX1 U1_4 (.A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]));
   FADDX1 U1_3 (.A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]));
   FADDX1 U1_2 (.A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]));
   FADDX1 U1_1 (.A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]));
   XOR3X1 U1_15 (.IN1(A[15]), .IN2(B[15]), .IN3(carry[15]), .Q(SUM[15]));
   AND2X1 U1 (.IN1(A[0]), .IN2(B[0]), .Q(n1));
   XOR2X1 U2 (.IN1(A[0]), .IN2(B[0]), .Q(SUM[0]));
endmodule

module ALU (a, b, alu_control, result, zero);
input [15:0] a;
input [15:0] b;
input [2:0] alu_control;
output zero;
output [15:0] result;
wire N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, 
       N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N79, N80
       , N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, 
       N97, N98, N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, 
       N143, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, 
       n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79
       , n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
       n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, 
       n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123
       , n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n1, n2, 
       n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n16, n17, n18, n19, n20, n21, n22, 
       n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
       , n40, n41, n42, n43, n44, n45, n46, n69, n136, n137, n138, n139, n140, n141, n142
       , n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n166, n167, 
       n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181
       , n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
       n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208
       , n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
       n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235
       , n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
       n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262
       , n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
       n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289
       , n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
       n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316
       , n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
       n330;
   NOR4X0 U56 (.IN1(n59), .IN2(n60), .IN3(n61), .IN4(n62), .QN(zero));
   OR4X1 U57 (.IN1(result[0]), .IN2(result[10]), .IN3(result[11]), .IN4(result[12]), .Q(
          n62));
   OR2X1 U58 (.IN1(n63), .IN2(n64), .Q(result[12]));
   AO222X1 U59 (.IN1(N59), .IN2(n65), .IN3(n66), .IN4(n178), .IN5(N43), .IN6(n67), .Q(n64)
          );
   AO221X1 U60 (.IN1(b[12]), .IN2(n68), .IN3(a[12]), .IN4(n9), .IN5(n70), .Q(n63));
   AO22X1 U61 (.IN1(N91), .IN2(n71), .IN3(N107), .IN4(n72), .Q(n70));
   AO21X1 U62 (.IN1(a[12]), .IN2(n73), .IN3(n10), .Q(n68));
   OR2X1 U63 (.IN1(n74), .IN2(n75), .Q(result[11]));
   AO222X1 U64 (.IN1(N58), .IN2(n65), .IN3(n66), .IN4(n181), .IN5(N42), .IN6(n67), .Q(n75)
          );
   AO221X1 U65 (.IN1(b[11]), .IN2(n76), .IN3(a[11]), .IN4(n9), .IN5(n77), .Q(n74));
   AO22X1 U66 (.IN1(N90), .IN2(n71), .IN3(N106), .IN4(n72), .Q(n77));
   AO21X1 U67 (.IN1(a[11]), .IN2(n73), .IN3(n10), .Q(n76));
   OR2X1 U68 (.IN1(n78), .IN2(n79), .Q(result[10]));
   AO222X1 U69 (.IN1(N57), .IN2(n65), .IN3(n66), .IN4(n186), .IN5(N41), .IN6(n67), .Q(n79)
          );
   AO221X1 U70 (.IN1(b[10]), .IN2(n80), .IN3(a[10]), .IN4(n9), .IN5(n81), .Q(n78));
   AO22X1 U71 (.IN1(N89), .IN2(n71), .IN3(N105), .IN4(n72), .Q(n81));
   AO21X1 U72 (.IN1(a[10]), .IN2(n73), .IN3(n9), .Q(n80));
   NAND4X0 U73 (.IN1(n82), .IN2(n83), .IN3(n84), .IN4(n85), .QN(result[0]));
   AOI221X1 U74 (.IN1(N79), .IN2(n71), .IN3(n66), .IN4(n206), .IN5(n86), .QN(n85));
   AO22X1 U75 (.IN1(N31), .IN2(n67), .IN3(N47), .IN4(n65), .Q(n86));
   AOI22X1 U76 (.IN1(a[0]), .IN2(n9), .IN3(N95), .IN4(n72), .QN(n84));
   NAND4X0 U77 (.IN1(N143), .IN2(alu_control[1]), .IN3(alu_control[2]), .IN4(
          alu_control[0]), .QN(n83));
   AO21X1 U78 (.IN1(a[0]), .IN2(n73), .IN3(n9), .Q(n87));
   NAND4X0 U79 (.IN1(n58), .IN2(n57), .IN3(n56), .IN4(n55), .QN(n61));
   AO222X1 U80 (.IN1(N48), .IN2(n65), .IN3(n66), .IN4(n204), .IN5(N32), .IN6(n67), .Q(n89)
          );
   AO221X1 U81 (.IN1(n6), .IN2(n90), .IN3(a[1]), .IN4(n9), .IN5(n91), .Q(n88));
   AO22X1 U82 (.IN1(N80), .IN2(n71), .IN3(N96), .IN4(n72), .Q(n91));
   AO21X1 U83 (.IN1(a[1]), .IN2(n73), .IN3(n10), .Q(n90));
   AO222X1 U84 (.IN1(N62), .IN2(n65), .IN3(n66), .IN4(n169), .IN5(N46), .IN6(n67), .Q(n93)
          );
   AO221X1 U85 (.IN1(b[15]), .IN2(n94), .IN3(a[15]), .IN4(n9), .IN5(n95), .Q(n92));
   AO22X1 U86 (.IN1(N94), .IN2(n71), .IN3(N110), .IN4(n72), .Q(n95));
   AO21X1 U87 (.IN1(a[15]), .IN2(n73), .IN3(n9), .Q(n94));
   AO222X1 U88 (.IN1(N61), .IN2(n65), .IN3(n66), .IN4(n173), .IN5(N45), .IN6(n67), .Q(n97)
          );
   AO221X1 U89 (.IN1(b[14]), .IN2(n98), .IN3(a[14]), .IN4(n9), .IN5(n99), .Q(n96));
   AO22X1 U90 (.IN1(N93), .IN2(n71), .IN3(N109), .IN4(n72), .Q(n99));
   AO21X1 U91 (.IN1(a[14]), .IN2(n73), .IN3(n10), .Q(n98));
   AO222X1 U92 (.IN1(N60), .IN2(n65), .IN3(n66), .IN4(n150), .IN5(N44), .IN6(n67), .Q(n101)
          );
   AO221X1 U93 (.IN1(b[13]), .IN2(n102), .IN3(a[13]), .IN4(n9), .IN5(n103), .Q(n100));
   AO22X1 U94 (.IN1(N92), .IN2(n71), .IN3(N108), .IN4(n72), .Q(n103));
   AO21X1 U95 (.IN1(a[13]), .IN2(n73), .IN3(n10), .Q(n102));
   NAND4X0 U96 (.IN1(n54), .IN2(n53), .IN3(n52), .IN4(n51), .QN(n60));
   AO222X1 U97 (.IN1(N52), .IN2(n65), .IN3(n66), .IN4(n142), .IN5(N36), .IN6(n67), .Q(n105)
          );
   AO221X1 U98 (.IN1(b[5]), .IN2(n106), .IN3(a[5]), .IN4(n9), .IN5(n107), .Q(n104));
   AO22X1 U99 (.IN1(N84), .IN2(n71), .IN3(N100), .IN4(n72), .Q(n107));
   AO21X1 U100 (.IN1(a[5]), .IN2(n73), .IN3(n10), .Q(n106));
   AO222X1 U101 (.IN1(N51), .IN2(n65), .IN3(n66), .IN4(n199), .IN5(N35), .IN6(n67), .Q(
          n109));
   AO221X1 U102 (.IN1(b[4]), .IN2(n110), .IN3(a[4]), .IN4(n10), .IN5(n111), .Q(n108));
   AO22X1 U103 (.IN1(N83), .IN2(n71), .IN3(N99), .IN4(n72), .Q(n111));
   AO21X1 U104 (.IN1(a[4]), .IN2(n73), .IN3(n10), .Q(n110));
   AO222X1 U105 (.IN1(N50), .IN2(n65), .IN3(n66), .IN4(n200), .IN5(N34), .IN6(n67), .Q(
          n113));
   AO221X1 U106 (.IN1(n2), .IN2(n114), .IN3(a[3]), .IN4(n9), .IN5(n115), .Q(n112));
   AO22X1 U107 (.IN1(N82), .IN2(n71), .IN3(N98), .IN4(n72), .Q(n115));
   AO21X1 U108 (.IN1(a[3]), .IN2(n73), .IN3(n10), .Q(n114));
   AO222X1 U109 (.IN1(N49), .IN2(n65), .IN3(n66), .IN4(n202), .IN5(N33), .IN6(n67), .Q(
          n117));
   AO221X1 U110 (.IN1(n8), .IN2(n118), .IN3(a[2]), .IN4(n10), .IN5(n119), .Q(n116));
   AO22X1 U111 (.IN1(N81), .IN2(n71), .IN3(N97), .IN4(n72), .Q(n119));
   AO21X1 U112 (.IN1(a[2]), .IN2(n73), .IN3(n10), .Q(n118));
   NAND4X0 U113 (.IN1(n50), .IN2(n49), .IN3(n48), .IN4(n47), .QN(n59));
   AO222X1 U114 (.IN1(N56), .IN2(n65), .IN3(n66), .IN4(n146), .IN5(N40), .IN6(n67), .Q(
          n121));
   AO221X1 U115 (.IN1(b[9]), .IN2(n122), .IN3(n10), .IN4(a[9]), .IN5(n123), .Q(n120));
   AO22X1 U116 (.IN1(N88), .IN2(n71), .IN3(N104), .IN4(n72), .Q(n123));
   AO21X1 U117 (.IN1(a[9]), .IN2(n73), .IN3(n10), .Q(n122));
   AO222X1 U118 (.IN1(N55), .IN2(n65), .IN3(n66), .IN4(n191), .IN5(N39), .IN6(n67), .Q(
          n125));
   AO221X1 U119 (.IN1(b[8]), .IN2(n126), .IN3(a[8]), .IN4(n9), .IN5(n127), .Q(n124));
   AO22X1 U120 (.IN1(N87), .IN2(n71), .IN3(N103), .IN4(n72), .Q(n127));
   AO21X1 U121 (.IN1(a[8]), .IN2(n73), .IN3(n10), .Q(n126));
   AO222X1 U122 (.IN1(N54), .IN2(n65), .IN3(n66), .IN4(n193), .IN5(N38), .IN6(n67), .Q(
          n129));
   AO221X1 U123 (.IN1(b[7]), .IN2(n130), .IN3(a[7]), .IN4(n9), .IN5(n131), .Q(n128));
   AO22X1 U124 (.IN1(N86), .IN2(n71), .IN3(N102), .IN4(n72), .Q(n131));
   AO21X1 U125 (.IN1(a[7]), .IN2(n73), .IN3(n10), .Q(n130));
   AO222X1 U126 (.IN1(N53), .IN2(n65), .IN3(n66), .IN4(n196), .IN5(N37), .IN6(n67), .Q(
          n133));
   NOR3X0 U127 (.IN1(alu_control[1]), .IN2(alu_control[2]), .IN3(alu_control[0]), .QN(n67)
          );
   NOR3X0 U128 (.IN1(alu_control[0]), .IN2(alu_control[2]), .IN3(n210), .QN(n66));
   NOR3X0 U129 (.IN1(alu_control[1]), .IN2(alu_control[2]), .IN3(n208), .QN(n65));
   AO221X1 U130 (.IN1(b[6]), .IN2(n134), .IN3(a[6]), .IN4(n9), .IN5(n135), .Q(n132));
   AO22X1 U131 (.IN1(N85), .IN2(n71), .IN3(N101), .IN4(n72), .Q(n135));
   NOR3X0 U132 (.IN1(alu_control[0]), .IN2(alu_control[1]), .IN3(n209), .QN(n72));
   NOR3X0 U133 (.IN1(n208), .IN2(alu_control[2]), .IN3(n210), .QN(n71));
   AO21X1 U134 (.IN1(a[6]), .IN2(n73), .IN3(n10), .Q(n134));
   NOR3X0 U136 (.IN1(n208), .IN2(alu_control[1]), .IN3(n209), .QN(n73));
   ALU_DW01_sub_0 sub_17 (.A(a), .B({b[15:3], n8, n6, n4}), .CI(1'b0), .DIFF({N62, N61, 
          N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47}));
   ALU_DW01_add_0_DW01_add_2 add_16 (.A(a), .B({b[15:4], n2, n7, n5, n3}), .CI(1'b0), .SUM(
          {N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31})
          );
   OR3X1 U2 (.IN1(n209), .IN2(alu_control[0]), .IN3(n210), .Q(n1));
   INVX0 U3 (.INP(b[4]), .ZN(n12));
   INVX0 U4 (.INP(b[3]), .ZN(n11));
   INVX0 U5 (.INP(n260), .ZN(n192));
   INVX0 U6 (.INP(n257), .ZN(n198));
   INVX0 U7 (.INP(n329), .ZN(n166));
   INVX0 U8 (.INP(n259), .ZN(n194));
   INVX0 U9 (.INP(n330), .ZN(n168));
   INVX0 U12 (.INP(n4), .ZN(n207));
   INVX0 U13 (.INP(n8), .ZN(n203));
   INVX0 U14 (.INP(n6), .ZN(n205));
   INVX0 U15 (.INP(n292), .ZN(n171));
   INVX0 U16 (.INP(n253), .ZN(n170));
   INVX0 U17 (.INP(n1), .ZN(n10));
   INVX0 U18 (.INP(n1), .ZN(n9));
   INVX0 U19 (.INP(n241), .ZN(n195));
   INVX0 U20 (.INP(n267), .ZN(n197));
   INVX0 U21 (.INP(n319), .ZN(n175));
   INVX0 U22 (.INP(n286), .ZN(n167));
   INVX0 U23 (.INP(n324), .ZN(n185));
   INVX0 U24 (.INP(n314), .ZN(n190));
   NAND2X1 U25 (.IN1(n286), .IN2(n203), .QN(n326));
   NAND2X1 U26 (.IN1(n250), .IN2(n203), .QN(n256));
   NAND2X1 U27 (.IN1(n283), .IN2(n203), .QN(n312));
   NAND2X1 U28 (.IN1(n225), .IN2(n203), .QN(n264));
   INVX0 U29 (.INP(n268), .ZN(n187));
   INVX0 U30 (.INP(n263), .ZN(n189));
   INVX0 U31 (.INP(n217), .ZN(n179));
   INVX0 U32 (.INP(n214), .ZN(n182));
   INVX0 U33 (.INP(n321), .ZN(n176));
   INVX0 U34 (.INP(n311), .ZN(n180));
   INVX2 U35 (.INP(n11), .ZN(n2));
   INVX0 U36 (.INP(n55), .ZN(result[1]));
   INVX0 U37 (.INP(n54), .ZN(result[2]));
   NBUFFX4 U38 (.INP(b[1]), .Z(n6));
   NBUFFX4 U39 (.INP(b[2]), .Z(n8));
   NBUFFX4 U40 (.INP(b[0]), .Z(n4));
   NBUFFX2 U41 (.INP(b[1]), .Z(n5));
   INVX0 U42 (.INP(alu_control[2]), .ZN(n209));
   NBUFFX2 U43 (.INP(b[2]), .Z(n7));
   NBUFFX2 U44 (.INP(b[0]), .Z(n3));
   NOR2X0 U45 (.IN1(n284), .IN2(n5), .QN(n286));
   NOR2X0 U46 (.IN1(n215), .IN2(n5), .QN(n225));
   INVX0 U47 (.INP(alu_control[0]), .ZN(n208));
   INVX0 U48 (.INP(b[8]), .ZN(n145));
   INVX0 U49 (.INP(b[12]), .ZN(n149));
   INVX0 U50 (.INP(n224), .ZN(n201));
   INVX0 U51 (.INP(n303), .ZN(n183));
   INVX0 U52 (.INP(b[7]), .ZN(n143));
   INVX0 U53 (.INP(b[15]), .ZN(n151));
   INVX0 U54 (.INP(b[11]), .ZN(n147));
   NAND2X1 U55 (.IN1(n280), .IN2(n205), .QN(n285));
   NAND2X1 U135 (.IN1(n233), .IN2(n205), .QN(n254));
   INVX0 U137 (.INP(n136), .ZN(n153));
   INVX0 U138 (.INP(n69), .ZN(n148));
   INVX0 U139 (.INP(n232), .ZN(n174));
   INVX0 U140 (.INP(n298), .ZN(n188));
   INVX0 U141 (.INP(n306), .ZN(n184));
   INVX0 U142 (.INP(n47), .ZN(result[9]));
   NOR2X0 U143 (.IN1(n88), .IN2(n89), .QN(n55));
   INVX0 U144 (.INP(n53), .ZN(result[3]));
   INVX0 U145 (.INP(n52), .ZN(result[4]));
   INVX0 U146 (.INP(n51), .ZN(result[5]));
   INVX0 U147 (.INP(n50), .ZN(result[6]));
   INVX0 U148 (.INP(n49), .ZN(result[7]));
   INVX0 U149 (.INP(n48), .ZN(result[8]));
   INVX0 U150 (.INP(n58), .ZN(result[13]));
   INVX0 U151 (.INP(n57), .ZN(result[14]));
   INVX0 U152 (.INP(n56), .ZN(result[15]));
   NOR2X0 U153 (.IN1(n116), .IN2(n117), .QN(n54));
   NAND2X1 U154 (.IN1(n3), .IN2(n87), .QN(n82));
   INVX0 U155 (.INP(a[0]), .ZN(n206));
   INVX0 U156 (.INP(alu_control[1]), .ZN(n210));
   INVX0 U157 (.INP(n40), .ZN(n152));
   NAND2X1 U158 (.IN1(a[15]), .IN2(n207), .QN(n284));
   NAND2X1 U159 (.IN1(a[0]), .IN2(n207), .QN(n215));
   INVX0 U160 (.INP(a[5]), .ZN(n142));
   INVX0 U161 (.INP(a[9]), .ZN(n146));
   INVX0 U162 (.INP(a[13]), .ZN(n150));
   NOR2X0 U163 (.IN1(n120), .IN2(n121), .QN(n47));
   NOR2X0 U164 (.IN1(n104), .IN2(n105), .QN(n51));
   INVX0 U165 (.INP(a[2]), .ZN(n202));
   NOR2X0 U166 (.IN1(n124), .IN2(n125), .QN(n48));
   INVX0 U167 (.INP(a[8]), .ZN(n191));
   NOR2X0 U168 (.IN1(n108), .IN2(n109), .QN(n52));
   INVX0 U169 (.INP(a[4]), .ZN(n199));
   NOR2X0 U170 (.IN1(n92), .IN2(n93), .QN(n56));
   NOR2X0 U171 (.IN1(n128), .IN2(n129), .QN(n49));
   INVX0 U172 (.INP(a[7]), .ZN(n193));
   NOR2X0 U173 (.IN1(n112), .IN2(n113), .QN(n53));
   INVX0 U174 (.INP(a[3]), .ZN(n200));
   NOR2X0 U175 (.IN1(n96), .IN2(n97), .QN(n57));
   INVX0 U176 (.INP(a[14]), .ZN(n173));
   NOR2X0 U177 (.IN1(n132), .IN2(n133), .QN(n50));
   INVX0 U178 (.INP(a[6]), .ZN(n196));
   NOR2X0 U179 (.IN1(n100), .IN2(n101), .QN(n58));
   INVX0 U180 (.INP(a[1]), .ZN(n204));
   INVX0 U181 (.INP(a[15]), .ZN(n169));
   INVX0 U182 (.INP(n17), .ZN(n144));
   INVX0 U183 (.INP(a[11]), .ZN(n181));
   INVX0 U184 (.INP(a[10]), .ZN(n186));
   INVX0 U185 (.INP(a[12]), .ZN(n178));
   INVX0 U186 (.INP(n281), .ZN(n177));
   INVX0 U187 (.INP(n282), .ZN(n172));
   NOR2X0 U188 (.IN1(n143), .IN2(a[7]), .QN(n13));
   AOI21X1 U189 (.IN1(b[6]), .IN2(n196), .IN3(n13), .QN(n28));
   NOR2X0 U190 (.IN1(b[6]), .IN2(n13), .QN(n16));
   AO22X1 U191 (.IN1(a[7]), .IN2(n143), .IN3(n16), .IN4(a[6]), .Q(n17));
   NOR2X0 U192 (.IN1(n28), .IN2(n17), .QN(n31));
   NAND2X0 U193 (.IN1(b[5]), .IN2(n142), .QN(n23));
   NAND2X0 U194 (.IN1(n23), .IN2(n12), .QN(n18));
   OA221X1 U195 (.IN1(n199), .IN2(n18), .IN3(b[5]), .IN4(n142), .IN5(n144), .Q(n30));
   NAND2X0 U196 (.IN1(n4), .IN2(n206), .QN(n21));
   OR2X1 U197 (.IN1(n205), .IN2(a[1]), .Q(n20));
   NOR2X0 U198 (.IN1(n11), .IN2(a[3]), .QN(n22));
   NOR2X0 U199 (.IN1(n8), .IN2(n22), .QN(n19));
   AO22X1 U200 (.IN1(a[3]), .IN2(n11), .IN3(n19), .IN4(a[2]), .Q(n24));
   AO221X1 U201 (.IN1(a[1]), .IN2(n205), .IN3(n21), .IN4(n20), .IN5(n24), .Q(n27));
   AOI21X1 U202 (.IN1(n202), .IN2(n8), .IN3(n22), .QN(n25));
   OA221X1 U203 (.IN1(n25), .IN2(n24), .IN3(a[4]), .IN4(n12), .IN5(n23), .Q(n26));
   NAND3X0 U204 (.IN1(n28), .IN2(n27), .IN3(n26), .QN(n29));
   OA21X1 U205 (.IN1(n31), .IN2(n30), .IN3(n29), .Q(n141));
   NAND2X0 U206 (.IN1(b[13]), .IN2(n150), .QN(n42));
   NAND3X0 U207 (.IN1(n42), .IN2(n149), .IN3(a[12]), .QN(n32));
   OA21X1 U208 (.IN1(b[13]), .IN2(n150), .IN3(n32), .Q(n36));
   NOR2X0 U209 (.IN1(n151), .IN2(a[15]), .QN(n34));
   NOR2X0 U210 (.IN1(b[14]), .IN2(n34), .QN(n33));
   AOI22X1 U211 (.IN1(a[15]), .IN2(n151), .IN3(n33), .IN4(a[14]), .QN(n35));
   AO21X1 U212 (.IN1(b[14]), .IN2(n173), .IN3(n34), .Q(n40));
   AO22X1 U213 (.IN1(n36), .IN2(n35), .IN3(n35), .IN4(n40), .Q(n46));
   NOR2X0 U214 (.IN1(n147), .IN2(a[11]), .QN(n38));
   NOR2X0 U215 (.IN1(b[10]), .IN2(n38), .QN(n37));
   AOI22X1 U216 (.IN1(a[11]), .IN2(n147), .IN3(n37), .IN4(a[10]), .QN(n44));
   AO21X1 U217 (.IN1(b[10]), .IN2(n186), .IN3(n38), .Q(n69));
   NAND2X0 U218 (.IN1(b[9]), .IN2(n146), .QN(n138));
   NAND3X0 U219 (.IN1(n138), .IN2(n145), .IN3(a[8]), .QN(n39));
   OA21X1 U220 (.IN1(b[9]), .IN2(n146), .IN3(n39), .Q(n43));
   OR2X1 U221 (.IN1(n149), .IN2(a[12]), .Q(n41));
   NAND3X0 U222 (.IN1(n42), .IN2(n41), .IN3(n152), .QN(n136));
   AO221X1 U223 (.IN1(n44), .IN2(n69), .IN3(n43), .IN4(n44), .IN5(n136), .Q(n45));
   AND2X1 U224 (.IN1(n46), .IN2(n45), .Q(n140));
   OR2X1 U225 (.IN1(n145), .IN2(a[8]), .Q(n137));
   NAND4X0 U226 (.IN1(n148), .IN2(n153), .IN3(n138), .IN4(n137), .QN(n139));
   AO22X1 U227 (.IN1(n141), .IN2(n140), .IN3(n140), .IN4(n139), .Q(N143));
   OR3X1 U228 (.IN1(b[14]), .IN2(b[13]), .IN3(b[12]), .Q(n213));
   OR3X1 U229 (.IN1(b[9]), .IN2(b[8]), .IN3(b[7]), .Q(n211));
   OR4X1 U230 (.IN1(b[6]), .IN2(b[5]), .IN3(b[15]), .IN4(n211), .Q(n212));
   NOR4X0 U231 (.IN1(b[11]), .IN2(b[10]), .IN3(n213), .IN4(n212), .QN(n253));
   NOR4X0 U232 (.IN1(b[4]), .IN2(n2), .IN3(n170), .IN4(n264), .QN(N79));
   MUX21X1 U233 (.IN1(a[3]), .IN2(a[4]), .S(n207), .Q(n223));
   MUX21X1 U234 (.IN1(a[5]), .IN2(a[6]), .S(n207), .Q(n220));
   MUX21X1 U235 (.IN1(n223), .IN2(n220), .S(n205), .Q(n241));
   MUX21X1 U236 (.IN1(a[7]), .IN2(a[8]), .S(n207), .Q(n219));
   MUX21X1 U237 (.IN1(a[9]), .IN2(a[10]), .S(n207), .Q(n221));
   MUX21X1 U238 (.IN1(n219), .IN2(n221), .S(n205), .Q(n240));
   MUX21X1 U239 (.IN1(n241), .IN2(n240), .S(n203), .Q(n214));
   MUX21X1 U240 (.IN1(a[1]), .IN2(a[2]), .S(n207), .Q(n224));
   MUX21X1 U241 (.IN1(n215), .IN2(n201), .S(n205), .Q(n242));
   OR2X1 U242 (.IN1(n242), .IN2(n8), .Q(n255));
   MUX21X1 U243 (.IN1(n182), .IN2(n255), .S(n2), .Q(n216));
   NOR3X0 U244 (.IN1(n216), .IN2(b[4]), .IN3(n170), .QN(N89));
   MUX21X1 U245 (.IN1(a[4]), .IN2(a[5]), .S(n207), .Q(n234));
   MUX21X1 U246 (.IN1(a[6]), .IN2(a[7]), .S(n207), .Q(n229));
   MUX21X1 U247 (.IN1(n234), .IN2(n229), .S(n205), .Q(n249));
   MUX21X1 U248 (.IN1(a[8]), .IN2(a[9]), .S(n207), .Q(n228));
   MUX21X1 U249 (.IN1(a[10]), .IN2(a[11]), .S(n207), .Q(n230));
   MUX21X1 U250 (.IN1(n228), .IN2(n230), .S(n205), .Q(n248));
   MUX21X1 U251 (.IN1(n249), .IN2(n248), .S(n203), .Q(n217));
   MUX21X1 U252 (.IN1(a[0]), .IN2(a[1]), .S(n207), .Q(n233));
   MUX21X1 U253 (.IN1(a[2]), .IN2(a[3]), .S(n207), .Q(n235));
   MUX21X1 U254 (.IN1(n233), .IN2(n235), .S(n205), .Q(n250));
   MUX21X1 U255 (.IN1(n179), .IN2(n256), .S(n2), .Q(n218));
   NOR3X0 U256 (.IN1(n218), .IN2(b[4]), .IN3(n170), .QN(N90));
   MUX21X1 U257 (.IN1(n220), .IN2(n219), .S(n205), .Q(n261));
   MUX21X1 U258 (.IN1(a[11]), .IN2(a[12]), .S(n207), .Q(n238));
   MUX21X1 U259 (.IN1(n221), .IN2(n238), .S(n205), .Q(n222));
   MUX21X1 U260 (.IN1(n261), .IN2(n222), .S(n203), .Q(n226));
   MUX21X1 U261 (.IN1(n224), .IN2(n223), .S(n205), .Q(n262));
   MUX21X1 U262 (.IN1(n225), .IN2(n262), .S(n203), .Q(n257));
   MUX21X1 U263 (.IN1(n226), .IN2(n257), .S(n2), .Q(n227));
   AND3X1 U264 (.IN1(n227), .IN2(n12), .IN3(n253), .Q(N91));
   MUX21X1 U265 (.IN1(n229), .IN2(n228), .S(n205), .Q(n266));
   MUX21X1 U266 (.IN1(a[12]), .IN2(a[13]), .S(n207), .Q(n246));
   MUX21X1 U267 (.IN1(n230), .IN2(n246), .S(n205), .Q(n231));
   MUX21X1 U268 (.IN1(n266), .IN2(n231), .S(n203), .Q(n232));
   MUX21X1 U269 (.IN1(n235), .IN2(n234), .S(n205), .Q(n267));
   MUX21X1 U270 (.IN1(n254), .IN2(n197), .S(n203), .Q(n258));
   MUX21X1 U271 (.IN1(n174), .IN2(n258), .S(n2), .Q(n236));
   NOR3X0 U272 (.IN1(n236), .IN2(b[4]), .IN3(n170), .QN(N92));
   MUX21X1 U273 (.IN1(a[13]), .IN2(a[14]), .S(n207), .Q(n237));
   MUX21X1 U274 (.IN1(n238), .IN2(n237), .S(n205), .Q(n239));
   MUX21X1 U275 (.IN1(n240), .IN2(n239), .S(n203), .Q(n243));
   MUX21X1 U276 (.IN1(n242), .IN2(n195), .S(n203), .Q(n259));
   MUX21X1 U277 (.IN1(n243), .IN2(n194), .S(n2), .Q(n244));
   AND3X1 U278 (.IN1(n253), .IN2(n12), .IN3(n244), .Q(N93));
   MUX21X1 U279 (.IN1(a[14]), .IN2(a[15]), .S(n207), .Q(n245));
   MUX21X1 U280 (.IN1(n246), .IN2(n245), .S(n205), .Q(n247));
   MUX21X1 U281 (.IN1(n248), .IN2(n247), .S(n203), .Q(n251));
   MUX21X1 U282 (.IN1(n250), .IN2(n249), .S(n203), .Q(n260));
   MUX21X1 U283 (.IN1(n251), .IN2(n260), .S(n2), .Q(n252));
   AND3X1 U284 (.IN1(n253), .IN2(n12), .IN3(n252), .Q(N94));
   OR2X1 U285 (.IN1(n254), .IN2(n8), .Q(n269));
   NOR4X0 U286 (.IN1(b[4]), .IN2(n2), .IN3(n170), .IN4(n269), .QN(N80));
   NOR4X0 U287 (.IN1(b[4]), .IN2(n2), .IN3(n170), .IN4(n255), .QN(N81));
   NOR4X0 U288 (.IN1(b[4]), .IN2(n2), .IN3(n170), .IN4(n256), .QN(N82));
   NOR4X0 U289 (.IN1(b[4]), .IN2(n2), .IN3(n198), .IN4(n170), .QN(N83));
   NOR4X0 U290 (.IN1(b[4]), .IN2(n2), .IN3(n258), .IN4(n170), .QN(N84));
   NOR4X0 U291 (.IN1(b[4]), .IN2(n2), .IN3(n259), .IN4(n170), .QN(N85));
   NOR4X0 U292 (.IN1(b[4]), .IN2(n2), .IN3(n192), .IN4(n170), .QN(N86));
   MUX21X1 U293 (.IN1(n262), .IN2(n261), .S(n203), .Q(n263));
   MUX21X1 U294 (.IN1(n189), .IN2(n264), .S(n2), .Q(n265));
   NOR3X0 U295 (.IN1(n265), .IN2(b[4]), .IN3(n170), .QN(N87));
   MUX21X1 U296 (.IN1(n267), .IN2(n266), .S(n203), .Q(n268));
   MUX21X1 U297 (.IN1(n187), .IN2(n269), .S(n2), .Q(n270));
   NOR3X0 U298 (.IN1(n270), .IN2(b[4]), .IN3(n170), .QN(N88));
   OR3X1 U299 (.IN1(b[14]), .IN2(b[13]), .IN3(b[12]), .Q(n273));
   OR3X1 U300 (.IN1(b[9]), .IN2(b[8]), .IN3(b[7]), .Q(n271));
   OR4X1 U301 (.IN1(b[6]), .IN2(b[5]), .IN3(b[15]), .IN4(n271), .Q(n272));
   NOR4X0 U302 (.IN1(b[11]), .IN2(b[10]), .IN3(n273), .IN4(n272), .QN(n292));
   MUX21X1 U303 (.IN1(a[0]), .IN2(a[1]), .S(n4), .Q(n274));
   MUX21X1 U304 (.IN1(a[2]), .IN2(a[3]), .S(n4), .Q(n294));
   MUX21X1 U305 (.IN1(n274), .IN2(n294), .S(n6), .Q(n275));
   MUX21X1 U306 (.IN1(a[4]), .IN2(a[5]), .S(n4), .Q(n293));
   MUX21X1 U307 (.IN1(a[6]), .IN2(a[7]), .S(n4), .Q(n296));
   MUX21X1 U308 (.IN1(n293), .IN2(n296), .S(n6), .Q(n310));
   MUX21X1 U309 (.IN1(n275), .IN2(n310), .S(n7), .Q(n276));
   MUX21X1 U310 (.IN1(a[8]), .IN2(a[9]), .S(n4), .Q(n295));
   MUX21X1 U311 (.IN1(a[10]), .IN2(a[11]), .S(n4), .Q(n279));
   MUX21X1 U312 (.IN1(n295), .IN2(n279), .S(n6), .Q(n309));
   MUX21X1 U313 (.IN1(a[12]), .IN2(a[13]), .S(n4), .Q(n278));
   MUX21X1 U314 (.IN1(a[14]), .IN2(a[15]), .S(n4), .Q(n280));
   MUX21X1 U315 (.IN1(n278), .IN2(n280), .S(n6), .Q(n283));
   MUX21X1 U316 (.IN1(n309), .IN2(n283), .S(n8), .Q(n329));
   MUX21X1 U317 (.IN1(n276), .IN2(n329), .S(n2), .Q(n277));
   AND3X1 U318 (.IN1(n292), .IN2(n12), .IN3(n277), .Q(N95));
   MUX21X1 U319 (.IN1(n279), .IN2(n278), .S(n6), .Q(n319));
   MUX21X1 U320 (.IN1(n175), .IN2(n285), .S(n8), .Q(n299));
   NOR4X0 U321 (.IN1(b[4]), .IN2(n2), .IN3(n299), .IN4(n171), .QN(N105));
   MUX21X1 U322 (.IN1(a[11]), .IN2(a[12]), .S(n4), .Q(n281));
   MUX21X1 U323 (.IN1(a[13]), .IN2(a[14]), .S(n4), .Q(n282));
   MUX21X1 U324 (.IN1(n177), .IN2(n172), .S(n6), .Q(n325));
   MUX21X1 U325 (.IN1(n325), .IN2(n167), .S(n8), .Q(n307));
   NOR4X0 U326 (.IN1(b[4]), .IN2(n2), .IN3(n307), .IN4(n171), .QN(N106));
   NOR4X0 U327 (.IN1(b[4]), .IN2(n2), .IN3(n171), .IN4(n312), .QN(N107));
   MUX21X1 U328 (.IN1(n172), .IN2(n284), .S(n6), .Q(n289));
   OR2X1 U329 (.IN1(n289), .IN2(n8), .Q(n316));
   NOR4X0 U330 (.IN1(b[4]), .IN2(n2), .IN3(n171), .IN4(n316), .QN(N108));
   OR2X1 U331 (.IN1(n285), .IN2(n8), .Q(n322));
   NOR4X0 U332 (.IN1(b[4]), .IN2(n2), .IN3(n171), .IN4(n322), .QN(N109));
   NOR4X0 U333 (.IN1(b[4]), .IN2(n2), .IN3(n171), .IN4(n326), .QN(N110));
   MUX21X1 U334 (.IN1(a[1]), .IN2(a[2]), .S(n4), .Q(n287));
   MUX21X1 U335 (.IN1(a[3]), .IN2(a[4]), .S(n4), .Q(n302));
   MUX21X1 U336 (.IN1(n287), .IN2(n302), .S(n6), .Q(n288));
   MUX21X1 U337 (.IN1(a[5]), .IN2(a[6]), .S(n4), .Q(n301));
   MUX21X1 U338 (.IN1(a[7]), .IN2(a[8]), .S(n4), .Q(n304));
   MUX21X1 U339 (.IN1(n301), .IN2(n304), .S(n6), .Q(n314));
   MUX21X1 U340 (.IN1(n288), .IN2(n314), .S(n8), .Q(n290));
   MUX21X1 U341 (.IN1(a[9]), .IN2(a[10]), .S(n4), .Q(n303));
   MUX21X1 U342 (.IN1(n183), .IN2(n177), .S(n6), .Q(n315));
   MUX21X1 U343 (.IN1(n315), .IN2(n289), .S(n8), .Q(n330));
   MUX21X1 U344 (.IN1(n290), .IN2(n168), .S(n2), .Q(n291));
   AND3X1 U345 (.IN1(n292), .IN2(n12), .IN3(n291), .Q(N96));
   MUX21X1 U346 (.IN1(n294), .IN2(n293), .S(n6), .Q(n297));
   MUX21X1 U347 (.IN1(n296), .IN2(n295), .S(n6), .Q(n320));
   MUX21X1 U348 (.IN1(n297), .IN2(n320), .S(n8), .Q(n298));
   MUX21X1 U349 (.IN1(n188), .IN2(n299), .S(n2), .Q(n300));
   NOR3X0 U350 (.IN1(n300), .IN2(b[4]), .IN3(n171), .QN(N97));
   MUX21X1 U351 (.IN1(n302), .IN2(n301), .S(n6), .Q(n305));
   MUX21X1 U352 (.IN1(n304), .IN2(n303), .S(n6), .Q(n324));
   MUX21X1 U353 (.IN1(n305), .IN2(n324), .S(n8), .Q(n306));
   MUX21X1 U354 (.IN1(n184), .IN2(n307), .S(n2), .Q(n308));
   NOR3X0 U355 (.IN1(n308), .IN2(b[4]), .IN3(n171), .QN(N98));
   MUX21X1 U356 (.IN1(n310), .IN2(n309), .S(n8), .Q(n311));
   MUX21X1 U357 (.IN1(n180), .IN2(n312), .S(n2), .Q(n313));
   NOR3X0 U358 (.IN1(n313), .IN2(b[4]), .IN3(n171), .QN(N99));
   MUX21X1 U359 (.IN1(n190), .IN2(n315), .S(n8), .Q(n317));
   MUX21X1 U360 (.IN1(n317), .IN2(n316), .S(n2), .Q(n318));
   NOR3X0 U361 (.IN1(n318), .IN2(b[4]), .IN3(n171), .QN(N100));
   MUX21X1 U362 (.IN1(n320), .IN2(n319), .S(n8), .Q(n321));
   MUX21X1 U363 (.IN1(n176), .IN2(n322), .S(n2), .Q(n323));
   NOR3X0 U364 (.IN1(n323), .IN2(b[4]), .IN3(n171), .QN(N101));
   MUX21X1 U365 (.IN1(n185), .IN2(n325), .S(n8), .Q(n327));
   MUX21X1 U366 (.IN1(n327), .IN2(n326), .S(n2), .Q(n328));
   NOR3X0 U367 (.IN1(n328), .IN2(b[4]), .IN3(n171), .QN(N102));
   NOR4X0 U368 (.IN1(b[4]), .IN2(n2), .IN3(n166), .IN4(n171), .QN(N103));
   NOR4X0 U369 (.IN1(b[4]), .IN2(n2), .IN3(n330), .IN4(n171), .QN(N104));
endmodule

module Data_Memory_test_1 (clk, mem_access_addr, mem_write_data, mem_write_en, mem_read, 
       mem_read_data, test_si2, test_si1, test_so2, test_so1, test_se);
input clk, mem_write_en, mem_read, test_si2, test_si1, test_se;
input [15:0] mem_access_addr;
input [15:0] mem_write_data;
output test_so2, test_so1;
output [15:0] mem_read_data;
wire N12, N13, N14, \memory[7][15] , \memory[7][14] , \memory[7][13] , \memory[7][12] , 
       \memory[7][11] , \memory[7][10] , \memory[7][9] , \memory[7][8] , \memory[7][7] , 
       \memory[7][6] , \memory[7][5] , \memory[7][4] , \memory[7][3] , \memory[7][2] , 
       \memory[7][1] , \memory[7][0] , \memory[6][15] , \memory[6][14] , \memory[6][13] , 
       \memory[6][12] , \memory[6][11] , \memory[6][10] , \memory[6][9] , \memory[6][8] , 
       \memory[6][7] , \memory[6][6] , \memory[6][5] , \memory[6][4] , \memory[6][3] , 
       \memory[6][2] , \memory[6][1] , \memory[6][0] , \memory[5][15] , \memory[5][14] , 
       \memory[5][13] , \memory[5][12] , \memory[5][11] , \memory[5][10] , \memory[5][9] 
       , \memory[5][8] , \memory[5][7] , \memory[5][6] , \memory[5][5] , \memory[5][4] , 
       \memory[5][3] , \memory[5][2] , \memory[5][1] , \memory[5][0] , \memory[4][15] , 
       \memory[4][14] , \memory[4][13] , \memory[4][12] , \memory[4][11] , \memory[4][10] 
       , \memory[4][9] , \memory[4][8] , \memory[4][7] , \memory[4][6] , \memory[4][5] , 
       \memory[4][4] , \memory[4][3] , \memory[4][2] , \memory[4][1] , \memory[4][0] , 
       \memory[3][15] , \memory[3][14] , \memory[3][13] , \memory[3][12] , \memory[3][11] 
       , \memory[3][10] , \memory[3][9] , \memory[3][8] , \memory[3][7] , \memory[3][6] , 
       \memory[3][5] , \memory[3][4] , \memory[3][3] , \memory[3][2] , \memory[3][1] , 
       \memory[3][0] , \memory[2][15] , \memory[2][14] , \memory[2][13] , \memory[2][12] 
       , \memory[2][11] , \memory[2][10] , \memory[2][9] , \memory[2][8] , \memory[2][7] 
       , \memory[2][6] , \memory[2][5] , \memory[2][4] , \memory[2][3] , \memory[2][2] , 
       \memory[2][1] , \memory[2][0] , \memory[1][15] , \memory[1][14] , \memory[1][13] , 
       \memory[1][12] , \memory[1][11] , \memory[1][10] , \memory[1][9] , \memory[1][8] , 
       \memory[1][7] , \memory[1][6] , \memory[1][5] , \memory[1][4] , \memory[1][3] , 
       \memory[1][2] , \memory[1][1] , \memory[1][0] , \memory[0][15] , \memory[0][14] , 
       \memory[0][13] , \memory[0][12] , \memory[0][11] , \memory[0][10] , \memory[0][9] 
       , \memory[0][8] , \memory[0][7] , \memory[0][6] , \memory[0][5] , \memory[0][4] , 
       \memory[0][3] , \memory[0][2] , \memory[0][1] , \memory[0][0] , N33, N34, N35, N36
       , N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, n140, n141, n142, 
       n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156
       , n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, 
       n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183
       , n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
       n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210
       , n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
       n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237
       , n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
       n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264
       , n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, 
       n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n278, n279, n280
       , n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
       n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307
       , n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
       n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334
       , n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
       n348, n349, n350, n351, n352, n353, n354, n355, n358, n359, n360, n361, n362, n363
       , n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
       n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390
       , n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
       n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417
       , n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
       n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444
       , n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, 
       n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471
       , n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483;
   assign N12 = mem_access_addr[0];
   assign N13 = mem_access_addr[1];
   assign N14 = mem_access_addr[2];
   assign test_so1 = \memory[5][10] ;
   SDFFX1 \memory_reg[7][15]  (.D(n277), .SI(n358), .SE(test_se), .CLK(clk), .Q(
          \memory[7][15] ), .QN(test_so2));
   SDFFX1 \memory_reg[7][14]  (.D(n276), .SI(n359), .SE(test_se), .CLK(clk), .Q(
          \memory[7][14] ), .QN(n358));
   SDFFX1 \memory_reg[7][13]  (.D(n275), .SI(n360), .SE(test_se), .CLK(clk), .Q(
          \memory[7][13] ), .QN(n359));
   SDFFX1 \memory_reg[7][12]  (.D(n274), .SI(n361), .SE(test_se), .CLK(clk), .Q(
          \memory[7][12] ), .QN(n360));
   SDFFX1 \memory_reg[7][11]  (.D(n273), .SI(n362), .SE(test_se), .CLK(clk), .Q(
          \memory[7][11] ), .QN(n361));
   SDFFX1 \memory_reg[7][10]  (.D(n272), .SI(n363), .SE(test_se), .CLK(clk), .Q(
          \memory[7][10] ), .QN(n362));
   SDFFX1 \memory_reg[7][9]  (.D(n271), .SI(n364), .SE(test_se), .CLK(clk), .Q(
          \memory[7][9] ), .QN(n363));
   SDFFX1 \memory_reg[7][8]  (.D(n270), .SI(n365), .SE(test_se), .CLK(clk), .Q(
          \memory[7][8] ), .QN(n364));
   SDFFX1 \memory_reg[7][7]  (.D(n269), .SI(n366), .SE(test_se), .CLK(clk), .Q(
          \memory[7][7] ), .QN(n365));
   SDFFX1 \memory_reg[7][6]  (.D(n268), .SI(n367), .SE(test_se), .CLK(clk), .Q(
          \memory[7][6] ), .QN(n366));
   SDFFX1 \memory_reg[7][5]  (.D(n267), .SI(n368), .SE(test_se), .CLK(clk), .Q(
          \memory[7][5] ), .QN(n367));
   SDFFX1 \memory_reg[7][4]  (.D(n266), .SI(n369), .SE(test_se), .CLK(clk), .Q(
          \memory[7][4] ), .QN(n368));
   SDFFX1 \memory_reg[7][3]  (.D(n265), .SI(n370), .SE(test_se), .CLK(clk), .Q(
          \memory[7][3] ), .QN(n369));
   SDFFX1 \memory_reg[7][2]  (.D(n264), .SI(n371), .SE(test_se), .CLK(clk), .Q(
          \memory[7][2] ), .QN(n370));
   SDFFX1 \memory_reg[7][1]  (.D(n263), .SI(n372), .SE(test_se), .CLK(clk), .Q(
          \memory[7][1] ), .QN(n371));
   SDFFX1 \memory_reg[7][0]  (.D(n262), .SI(n373), .SE(test_se), .CLK(clk), .Q(
          \memory[7][0] ), .QN(n372));
   SDFFX1 \memory_reg[6][15]  (.D(n261), .SI(n374), .SE(test_se), .CLK(clk), .Q(
          \memory[6][15] ), .QN(n373));
   SDFFX1 \memory_reg[6][14]  (.D(n260), .SI(n375), .SE(test_se), .CLK(clk), .Q(
          \memory[6][14] ), .QN(n374));
   SDFFX1 \memory_reg[6][13]  (.D(n259), .SI(n376), .SE(test_se), .CLK(clk), .Q(
          \memory[6][13] ), .QN(n375));
   SDFFX1 \memory_reg[6][12]  (.D(n258), .SI(n377), .SE(test_se), .CLK(clk), .Q(
          \memory[6][12] ), .QN(n376));
   SDFFX1 \memory_reg[6][11]  (.D(n257), .SI(n378), .SE(test_se), .CLK(clk), .Q(
          \memory[6][11] ), .QN(n377));
   SDFFX1 \memory_reg[6][10]  (.D(n256), .SI(n379), .SE(test_se), .CLK(clk), .Q(
          \memory[6][10] ), .QN(n378));
   SDFFX1 \memory_reg[6][9]  (.D(n255), .SI(n380), .SE(test_se), .CLK(clk), .Q(
          \memory[6][9] ), .QN(n379));
   SDFFX1 \memory_reg[6][8]  (.D(n254), .SI(n381), .SE(test_se), .CLK(clk), .Q(
          \memory[6][8] ), .QN(n380));
   SDFFX1 \memory_reg[6][7]  (.D(n253), .SI(n382), .SE(test_se), .CLK(clk), .Q(
          \memory[6][7] ), .QN(n381));
   SDFFX1 \memory_reg[6][6]  (.D(n252), .SI(n383), .SE(test_se), .CLK(clk), .Q(
          \memory[6][6] ), .QN(n382));
   SDFFX1 \memory_reg[6][5]  (.D(n251), .SI(n384), .SE(test_se), .CLK(clk), .Q(
          \memory[6][5] ), .QN(n383));
   SDFFX1 \memory_reg[6][4]  (.D(n250), .SI(n385), .SE(test_se), .CLK(clk), .Q(
          \memory[6][4] ), .QN(n384));
   SDFFX1 \memory_reg[6][3]  (.D(n249), .SI(n386), .SE(test_se), .CLK(clk), .Q(
          \memory[6][3] ), .QN(n385));
   SDFFX1 \memory_reg[6][2]  (.D(n248), .SI(n387), .SE(test_se), .CLK(clk), .Q(
          \memory[6][2] ), .QN(n386));
   SDFFX1 \memory_reg[6][1]  (.D(n247), .SI(n388), .SE(test_se), .CLK(clk), .Q(
          \memory[6][1] ), .QN(n387));
   SDFFX1 \memory_reg[6][0]  (.D(n246), .SI(n389), .SE(test_se), .CLK(clk), .Q(
          \memory[6][0] ), .QN(n388));
   SDFFX1 \memory_reg[5][15]  (.D(n245), .SI(n390), .SE(test_se), .CLK(clk), .Q(
          \memory[5][15] ), .QN(n389));
   SDFFX1 \memory_reg[5][14]  (.D(n244), .SI(n391), .SE(test_se), .CLK(clk), .Q(
          \memory[5][14] ), .QN(n390));
   SDFFX1 \memory_reg[5][13]  (.D(n243), .SI(n392), .SE(test_se), .CLK(clk), .Q(
          \memory[5][13] ), .QN(n391));
   SDFFX1 \memory_reg[5][12]  (.D(n242), .SI(n393), .SE(test_se), .CLK(clk), .Q(
          \memory[5][12] ), .QN(n392));
   SDFFX1 \memory_reg[5][11]  (.D(n241), .SI(test_si2), .SE(test_se), .CLK(clk), .Q(
          \memory[5][11] ), .QN(n393));
   SDFFX1 \memory_reg[5][10]  (.D(n240), .SI(n394), .SE(test_se), .CLK(clk), .Q(
          \memory[5][10] ));
   SDFFX1 \memory_reg[5][9]  (.D(n239), .SI(n395), .SE(test_se), .CLK(clk), .Q(
          \memory[5][9] ), .QN(n394));
   SDFFX1 \memory_reg[5][8]  (.D(n238), .SI(n396), .SE(test_se), .CLK(clk), .Q(
          \memory[5][8] ), .QN(n395));
   SDFFX1 \memory_reg[5][7]  (.D(n237), .SI(n397), .SE(test_se), .CLK(clk), .Q(
          \memory[5][7] ), .QN(n396));
   SDFFX1 \memory_reg[5][6]  (.D(n236), .SI(n398), .SE(test_se), .CLK(clk), .Q(
          \memory[5][6] ), .QN(n397));
   SDFFX1 \memory_reg[5][5]  (.D(n235), .SI(n399), .SE(test_se), .CLK(clk), .Q(
          \memory[5][5] ), .QN(n398));
   SDFFX1 \memory_reg[5][4]  (.D(n234), .SI(n400), .SE(test_se), .CLK(clk), .Q(
          \memory[5][4] ), .QN(n399));
   SDFFX1 \memory_reg[5][3]  (.D(n233), .SI(n401), .SE(test_se), .CLK(clk), .Q(
          \memory[5][3] ), .QN(n400));
   SDFFX1 \memory_reg[5][2]  (.D(n232), .SI(n402), .SE(test_se), .CLK(clk), .Q(
          \memory[5][2] ), .QN(n401));
   SDFFX1 \memory_reg[5][1]  (.D(n231), .SI(n403), .SE(test_se), .CLK(clk), .Q(
          \memory[5][1] ), .QN(n402));
   SDFFX1 \memory_reg[5][0]  (.D(n230), .SI(n404), .SE(test_se), .CLK(clk), .Q(
          \memory[5][0] ), .QN(n403));
   SDFFX1 \memory_reg[4][15]  (.D(n229), .SI(n405), .SE(test_se), .CLK(clk), .Q(
          \memory[4][15] ), .QN(n404));
   SDFFX1 \memory_reg[4][14]  (.D(n228), .SI(n406), .SE(test_se), .CLK(clk), .Q(
          \memory[4][14] ), .QN(n405));
   SDFFX1 \memory_reg[4][13]  (.D(n227), .SI(n407), .SE(test_se), .CLK(clk), .Q(
          \memory[4][13] ), .QN(n406));
   SDFFX1 \memory_reg[4][12]  (.D(n226), .SI(n408), .SE(test_se), .CLK(clk), .Q(
          \memory[4][12] ), .QN(n407));
   SDFFX1 \memory_reg[4][11]  (.D(n225), .SI(n409), .SE(test_se), .CLK(clk), .Q(
          \memory[4][11] ), .QN(n408));
   SDFFX1 \memory_reg[4][10]  (.D(n224), .SI(n410), .SE(test_se), .CLK(clk), .Q(
          \memory[4][10] ), .QN(n409));
   SDFFX1 \memory_reg[4][9]  (.D(n223), .SI(n411), .SE(test_se), .CLK(clk), .Q(
          \memory[4][9] ), .QN(n410));
   SDFFX1 \memory_reg[4][8]  (.D(n222), .SI(n412), .SE(test_se), .CLK(clk), .Q(
          \memory[4][8] ), .QN(n411));
   SDFFX1 \memory_reg[4][7]  (.D(n221), .SI(n413), .SE(test_se), .CLK(clk), .Q(
          \memory[4][7] ), .QN(n412));
   SDFFX1 \memory_reg[4][6]  (.D(n220), .SI(n414), .SE(test_se), .CLK(clk), .Q(
          \memory[4][6] ), .QN(n413));
   SDFFX1 \memory_reg[4][5]  (.D(n219), .SI(n415), .SE(test_se), .CLK(clk), .Q(
          \memory[4][5] ), .QN(n414));
   SDFFX1 \memory_reg[4][4]  (.D(n218), .SI(n416), .SE(test_se), .CLK(clk), .Q(
          \memory[4][4] ), .QN(n415));
   SDFFX1 \memory_reg[4][3]  (.D(n217), .SI(n417), .SE(test_se), .CLK(clk), .Q(
          \memory[4][3] ), .QN(n416));
   SDFFX1 \memory_reg[4][2]  (.D(n216), .SI(n418), .SE(test_se), .CLK(clk), .Q(
          \memory[4][2] ), .QN(n417));
   SDFFX1 \memory_reg[4][1]  (.D(n215), .SI(n419), .SE(test_se), .CLK(clk), .Q(
          \memory[4][1] ), .QN(n418));
   SDFFX1 \memory_reg[4][0]  (.D(n214), .SI(n420), .SE(test_se), .CLK(clk), .Q(
          \memory[4][0] ), .QN(n419));
   SDFFX1 \memory_reg[3][15]  (.D(n213), .SI(n421), .SE(test_se), .CLK(clk), .Q(
          \memory[3][15] ), .QN(n420));
   SDFFX1 \memory_reg[3][14]  (.D(n212), .SI(n422), .SE(test_se), .CLK(clk), .Q(
          \memory[3][14] ), .QN(n421));
   SDFFX1 \memory_reg[3][13]  (.D(n211), .SI(n423), .SE(test_se), .CLK(clk), .Q(
          \memory[3][13] ), .QN(n422));
   SDFFX1 \memory_reg[3][12]  (.D(n210), .SI(n424), .SE(test_se), .CLK(clk), .Q(
          \memory[3][12] ), .QN(n423));
   SDFFX1 \memory_reg[3][11]  (.D(n209), .SI(n425), .SE(test_se), .CLK(clk), .Q(
          \memory[3][11] ), .QN(n424));
   SDFFX1 \memory_reg[3][10]  (.D(n208), .SI(n426), .SE(test_se), .CLK(clk), .Q(
          \memory[3][10] ), .QN(n425));
   SDFFX1 \memory_reg[3][9]  (.D(n207), .SI(n427), .SE(test_se), .CLK(clk), .Q(
          \memory[3][9] ), .QN(n426));
   SDFFX1 \memory_reg[3][8]  (.D(n206), .SI(n428), .SE(test_se), .CLK(clk), .Q(
          \memory[3][8] ), .QN(n427));
   SDFFX1 \memory_reg[3][7]  (.D(n205), .SI(n429), .SE(test_se), .CLK(clk), .Q(
          \memory[3][7] ), .QN(n428));
   SDFFX1 \memory_reg[3][6]  (.D(n204), .SI(n430), .SE(test_se), .CLK(clk), .Q(
          \memory[3][6] ), .QN(n429));
   SDFFX1 \memory_reg[3][5]  (.D(n203), .SI(n431), .SE(test_se), .CLK(clk), .Q(
          \memory[3][5] ), .QN(n430));
   SDFFX1 \memory_reg[3][4]  (.D(n202), .SI(n432), .SE(test_se), .CLK(clk), .Q(
          \memory[3][4] ), .QN(n431));
   SDFFX1 \memory_reg[3][3]  (.D(n201), .SI(n433), .SE(test_se), .CLK(clk), .Q(
          \memory[3][3] ), .QN(n432));
   SDFFX1 \memory_reg[3][2]  (.D(n200), .SI(n434), .SE(test_se), .CLK(clk), .Q(
          \memory[3][2] ), .QN(n433));
   SDFFX1 \memory_reg[3][1]  (.D(n199), .SI(n435), .SE(test_se), .CLK(clk), .Q(
          \memory[3][1] ), .QN(n434));
   SDFFX1 \memory_reg[3][0]  (.D(n198), .SI(n436), .SE(test_se), .CLK(clk), .Q(
          \memory[3][0] ), .QN(n435));
   SDFFX1 \memory_reg[2][15]  (.D(n197), .SI(n437), .SE(test_se), .CLK(clk), .Q(
          \memory[2][15] ), .QN(n436));
   SDFFX1 \memory_reg[2][14]  (.D(n196), .SI(n438), .SE(test_se), .CLK(clk), .Q(
          \memory[2][14] ), .QN(n437));
   SDFFX1 \memory_reg[2][13]  (.D(n195), .SI(n439), .SE(test_se), .CLK(clk), .Q(
          \memory[2][13] ), .QN(n438));
   SDFFX1 \memory_reg[2][12]  (.D(n194), .SI(n440), .SE(test_se), .CLK(clk), .Q(
          \memory[2][12] ), .QN(n439));
   SDFFX1 \memory_reg[2][11]  (.D(n193), .SI(n441), .SE(test_se), .CLK(clk), .Q(
          \memory[2][11] ), .QN(n440));
   SDFFX1 \memory_reg[2][10]  (.D(n192), .SI(n442), .SE(test_se), .CLK(clk), .Q(
          \memory[2][10] ), .QN(n441));
   SDFFX1 \memory_reg[2][9]  (.D(n191), .SI(n443), .SE(test_se), .CLK(clk), .Q(
          \memory[2][9] ), .QN(n442));
   SDFFX1 \memory_reg[2][8]  (.D(n190), .SI(n444), .SE(test_se), .CLK(clk), .Q(
          \memory[2][8] ), .QN(n443));
   SDFFX1 \memory_reg[2][7]  (.D(n189), .SI(n445), .SE(test_se), .CLK(clk), .Q(
          \memory[2][7] ), .QN(n444));
   SDFFX1 \memory_reg[2][6]  (.D(n188), .SI(n446), .SE(test_se), .CLK(clk), .Q(
          \memory[2][6] ), .QN(n445));
   SDFFX1 \memory_reg[2][5]  (.D(n187), .SI(n447), .SE(test_se), .CLK(clk), .Q(
          \memory[2][5] ), .QN(n446));
   SDFFX1 \memory_reg[2][4]  (.D(n186), .SI(n448), .SE(test_se), .CLK(clk), .Q(
          \memory[2][4] ), .QN(n447));
   SDFFX1 \memory_reg[2][3]  (.D(n185), .SI(n449), .SE(test_se), .CLK(clk), .Q(
          \memory[2][3] ), .QN(n448));
   SDFFX1 \memory_reg[2][2]  (.D(n184), .SI(n450), .SE(test_se), .CLK(clk), .Q(
          \memory[2][2] ), .QN(n449));
   SDFFX1 \memory_reg[2][1]  (.D(n183), .SI(n451), .SE(test_se), .CLK(clk), .Q(
          \memory[2][1] ), .QN(n450));
   SDFFX1 \memory_reg[2][0]  (.D(n182), .SI(n452), .SE(test_se), .CLK(clk), .Q(
          \memory[2][0] ), .QN(n451));
   SDFFX1 \memory_reg[1][15]  (.D(n181), .SI(n453), .SE(test_se), .CLK(clk), .Q(
          \memory[1][15] ), .QN(n452));
   SDFFX1 \memory_reg[1][14]  (.D(n180), .SI(n454), .SE(test_se), .CLK(clk), .Q(
          \memory[1][14] ), .QN(n453));
   SDFFX1 \memory_reg[1][13]  (.D(n179), .SI(n455), .SE(test_se), .CLK(clk), .Q(
          \memory[1][13] ), .QN(n454));
   SDFFX1 \memory_reg[1][12]  (.D(n178), .SI(n456), .SE(test_se), .CLK(clk), .Q(
          \memory[1][12] ), .QN(n455));
   SDFFX1 \memory_reg[1][11]  (.D(n177), .SI(n457), .SE(test_se), .CLK(clk), .Q(
          \memory[1][11] ), .QN(n456));
   SDFFX1 \memory_reg[1][10]  (.D(n176), .SI(n458), .SE(test_se), .CLK(clk), .Q(
          \memory[1][10] ), .QN(n457));
   SDFFX1 \memory_reg[1][9]  (.D(n175), .SI(n459), .SE(test_se), .CLK(clk), .Q(
          \memory[1][9] ), .QN(n458));
   SDFFX1 \memory_reg[1][8]  (.D(n174), .SI(n460), .SE(test_se), .CLK(clk), .Q(
          \memory[1][8] ), .QN(n459));
   SDFFX1 \memory_reg[1][7]  (.D(n173), .SI(n461), .SE(test_se), .CLK(clk), .Q(
          \memory[1][7] ), .QN(n460));
   SDFFX1 \memory_reg[1][6]  (.D(n172), .SI(n462), .SE(test_se), .CLK(clk), .Q(
          \memory[1][6] ), .QN(n461));
   SDFFX1 \memory_reg[1][5]  (.D(n171), .SI(n463), .SE(test_se), .CLK(clk), .Q(
          \memory[1][5] ), .QN(n462));
   SDFFX1 \memory_reg[1][4]  (.D(n170), .SI(n464), .SE(test_se), .CLK(clk), .Q(
          \memory[1][4] ), .QN(n463));
   SDFFX1 \memory_reg[1][3]  (.D(n169), .SI(n465), .SE(test_se), .CLK(clk), .Q(
          \memory[1][3] ), .QN(n464));
   SDFFX1 \memory_reg[1][2]  (.D(n168), .SI(n466), .SE(test_se), .CLK(clk), .Q(
          \memory[1][2] ), .QN(n465));
   SDFFX1 \memory_reg[1][1]  (.D(n167), .SI(n467), .SE(test_se), .CLK(clk), .Q(
          \memory[1][1] ), .QN(n466));
   SDFFX1 \memory_reg[1][0]  (.D(n166), .SI(n468), .SE(test_se), .CLK(clk), .Q(
          \memory[1][0] ), .QN(n467));
   SDFFX1 \memory_reg[0][15]  (.D(n165), .SI(n469), .SE(test_se), .CLK(clk), .Q(
          \memory[0][15] ), .QN(n468));
   SDFFX1 \memory_reg[0][14]  (.D(n164), .SI(n470), .SE(test_se), .CLK(clk), .Q(
          \memory[0][14] ), .QN(n469));
   SDFFX1 \memory_reg[0][13]  (.D(n163), .SI(n471), .SE(test_se), .CLK(clk), .Q(
          \memory[0][13] ), .QN(n470));
   SDFFX1 \memory_reg[0][12]  (.D(n162), .SI(n472), .SE(test_se), .CLK(clk), .Q(
          \memory[0][12] ), .QN(n471));
   SDFFX1 \memory_reg[0][11]  (.D(n161), .SI(n473), .SE(test_se), .CLK(clk), .Q(
          \memory[0][11] ), .QN(n472));
   SDFFX1 \memory_reg[0][10]  (.D(n160), .SI(n474), .SE(test_se), .CLK(clk), .Q(
          \memory[0][10] ), .QN(n473));
   SDFFX1 \memory_reg[0][9]  (.D(n159), .SI(n475), .SE(test_se), .CLK(clk), .Q(
          \memory[0][9] ), .QN(n474));
   SDFFX1 \memory_reg[0][8]  (.D(n158), .SI(n476), .SE(test_se), .CLK(clk), .Q(
          \memory[0][8] ), .QN(n475));
   SDFFX1 \memory_reg[0][7]  (.D(n157), .SI(n477), .SE(test_se), .CLK(clk), .Q(
          \memory[0][7] ), .QN(n476));
   SDFFX1 \memory_reg[0][6]  (.D(n156), .SI(n478), .SE(test_se), .CLK(clk), .Q(
          \memory[0][6] ), .QN(n477));
   SDFFX1 \memory_reg[0][5]  (.D(n155), .SI(n479), .SE(test_se), .CLK(clk), .Q(
          \memory[0][5] ), .QN(n478));
   SDFFX1 \memory_reg[0][4]  (.D(n154), .SI(n480), .SE(test_se), .CLK(clk), .Q(
          \memory[0][4] ), .QN(n479));
   SDFFX1 \memory_reg[0][3]  (.D(n153), .SI(n481), .SE(test_se), .CLK(clk), .Q(
          \memory[0][3] ), .QN(n480));
   SDFFX1 \memory_reg[0][2]  (.D(n152), .SI(n482), .SE(test_se), .CLK(clk), .Q(
          \memory[0][2] ), .QN(n481));
   SDFFX1 \memory_reg[0][1]  (.D(n151), .SI(n483), .SE(test_se), .CLK(clk), .Q(
          \memory[0][1] ), .QN(n482));
   SDFFX1 \memory_reg[0][0]  (.D(n150), .SI(test_si1), .SE(test_se), .CLK(clk), .Q(
          \memory[0][0] ), .QN(n483));
   AO22X1 U142 (.IN1(mem_write_data[0]), .IN2(n349), .IN3(\memory[0][0] ), .IN4(n140), .Q(
          n150));
   AO22X1 U143 (.IN1(mem_write_data[1]), .IN2(n349), .IN3(\memory[0][1] ), .IN4(n140), .Q(
          n151));
   AO22X1 U144 (.IN1(mem_write_data[2]), .IN2(n349), .IN3(\memory[0][2] ), .IN4(n140), .Q(
          n152));
   AO22X1 U145 (.IN1(mem_write_data[3]), .IN2(n349), .IN3(\memory[0][3] ), .IN4(n140), .Q(
          n153));
   AO22X1 U146 (.IN1(mem_write_data[4]), .IN2(n349), .IN3(\memory[0][4] ), .IN4(n140), .Q(
          n154));
   AO22X1 U147 (.IN1(mem_write_data[5]), .IN2(n349), .IN3(\memory[0][5] ), .IN4(n140), .Q(
          n155));
   AO22X1 U148 (.IN1(mem_write_data[6]), .IN2(n349), .IN3(\memory[0][6] ), .IN4(n140), .Q(
          n156));
   AO22X1 U149 (.IN1(mem_write_data[7]), .IN2(n349), .IN3(\memory[0][7] ), .IN4(n140), .Q(
          n157));
   AO22X1 U150 (.IN1(mem_write_data[8]), .IN2(n349), .IN3(\memory[0][8] ), .IN4(n140), .Q(
          n158));
   AO22X1 U151 (.IN1(mem_write_data[9]), .IN2(n349), .IN3(\memory[0][9] ), .IN4(n140), .Q(
          n159));
   AO22X1 U152 (.IN1(mem_write_data[10]), .IN2(n349), .IN3(\memory[0][10] ), .IN4(n140), .
          Q(n160));
   AO22X1 U153 (.IN1(mem_write_data[11]), .IN2(n349), .IN3(\memory[0][11] ), .IN4(n140), .
          Q(n161));
   AO22X1 U154 (.IN1(mem_write_data[12]), .IN2(n349), .IN3(\memory[0][12] ), .IN4(n140), .
          Q(n162));
   AO22X1 U155 (.IN1(mem_write_data[13]), .IN2(n349), .IN3(\memory[0][13] ), .IN4(n140), .
          Q(n163));
   AO22X1 U156 (.IN1(mem_write_data[14]), .IN2(n349), .IN3(\memory[0][14] ), .IN4(n140), .
          Q(n164));
   AO22X1 U157 (.IN1(mem_write_data[15]), .IN2(n349), .IN3(\memory[0][15] ), .IN4(n140), .
          Q(n165));
   AO22X1 U159 (.IN1(n348), .IN2(mem_write_data[0]), .IN3(\memory[1][0] ), .IN4(n142), .Q(
          n166));
   AO22X1 U160 (.IN1(n348), .IN2(mem_write_data[1]), .IN3(\memory[1][1] ), .IN4(n142), .Q(
          n167));
   AO22X1 U161 (.IN1(n348), .IN2(mem_write_data[2]), .IN3(\memory[1][2] ), .IN4(n142), .Q(
          n168));
   AO22X1 U162 (.IN1(n348), .IN2(mem_write_data[3]), .IN3(\memory[1][3] ), .IN4(n142), .Q(
          n169));
   AO22X1 U163 (.IN1(n348), .IN2(mem_write_data[4]), .IN3(\memory[1][4] ), .IN4(n142), .Q(
          n170));
   AO22X1 U164 (.IN1(n348), .IN2(mem_write_data[5]), .IN3(\memory[1][5] ), .IN4(n142), .Q(
          n171));
   AO22X1 U165 (.IN1(n348), .IN2(mem_write_data[6]), .IN3(\memory[1][6] ), .IN4(n142), .Q(
          n172));
   AO22X1 U166 (.IN1(n348), .IN2(mem_write_data[7]), .IN3(\memory[1][7] ), .IN4(n142), .Q(
          n173));
   AO22X1 U167 (.IN1(n348), .IN2(mem_write_data[8]), .IN3(\memory[1][8] ), .IN4(n142), .Q(
          n174));
   AO22X1 U168 (.IN1(n348), .IN2(mem_write_data[9]), .IN3(\memory[1][9] ), .IN4(n142), .Q(
          n175));
   AO22X1 U169 (.IN1(n348), .IN2(mem_write_data[10]), .IN3(\memory[1][10] ), .IN4(n142), .
          Q(n176));
   AO22X1 U170 (.IN1(n348), .IN2(mem_write_data[11]), .IN3(\memory[1][11] ), .IN4(n142), .
          Q(n177));
   AO22X1 U171 (.IN1(n348), .IN2(mem_write_data[12]), .IN3(\memory[1][12] ), .IN4(n142), .
          Q(n178));
   AO22X1 U172 (.IN1(n348), .IN2(mem_write_data[13]), .IN3(\memory[1][13] ), .IN4(n142), .
          Q(n179));
   AO22X1 U173 (.IN1(n348), .IN2(mem_write_data[14]), .IN3(\memory[1][14] ), .IN4(n142), .
          Q(n180));
   AO22X1 U174 (.IN1(n348), .IN2(mem_write_data[15]), .IN3(\memory[1][15] ), .IN4(n142), .
          Q(n181));
   AO22X1 U176 (.IN1(n347), .IN2(mem_write_data[0]), .IN3(\memory[2][0] ), .IN4(n143), .Q(
          n182));
   AO22X1 U177 (.IN1(n347), .IN2(mem_write_data[1]), .IN3(\memory[2][1] ), .IN4(n143), .Q(
          n183));
   AO22X1 U178 (.IN1(n347), .IN2(mem_write_data[2]), .IN3(\memory[2][2] ), .IN4(n143), .Q(
          n184));
   AO22X1 U179 (.IN1(n347), .IN2(mem_write_data[3]), .IN3(\memory[2][3] ), .IN4(n143), .Q(
          n185));
   AO22X1 U180 (.IN1(n347), .IN2(mem_write_data[4]), .IN3(\memory[2][4] ), .IN4(n143), .Q(
          n186));
   AO22X1 U181 (.IN1(n347), .IN2(mem_write_data[5]), .IN3(\memory[2][5] ), .IN4(n143), .Q(
          n187));
   AO22X1 U182 (.IN1(n347), .IN2(mem_write_data[6]), .IN3(\memory[2][6] ), .IN4(n143), .Q(
          n188));
   AO22X1 U183 (.IN1(n347), .IN2(mem_write_data[7]), .IN3(\memory[2][7] ), .IN4(n143), .Q(
          n189));
   AO22X1 U184 (.IN1(n347), .IN2(mem_write_data[8]), .IN3(\memory[2][8] ), .IN4(n143), .Q(
          n190));
   AO22X1 U185 (.IN1(n347), .IN2(mem_write_data[9]), .IN3(\memory[2][9] ), .IN4(n143), .Q(
          n191));
   AO22X1 U186 (.IN1(n347), .IN2(mem_write_data[10]), .IN3(\memory[2][10] ), .IN4(n143), .
          Q(n192));
   AO22X1 U187 (.IN1(n347), .IN2(mem_write_data[11]), .IN3(\memory[2][11] ), .IN4(n143), .
          Q(n193));
   AO22X1 U188 (.IN1(n347), .IN2(mem_write_data[12]), .IN3(\memory[2][12] ), .IN4(n143), .
          Q(n194));
   AO22X1 U189 (.IN1(n347), .IN2(mem_write_data[13]), .IN3(\memory[2][13] ), .IN4(n143), .
          Q(n195));
   AO22X1 U190 (.IN1(n347), .IN2(mem_write_data[14]), .IN3(\memory[2][14] ), .IN4(n143), .
          Q(n196));
   AO22X1 U191 (.IN1(n347), .IN2(mem_write_data[15]), .IN3(\memory[2][15] ), .IN4(n143), .
          Q(n197));
   AO22X1 U193 (.IN1(n346), .IN2(mem_write_data[0]), .IN3(\memory[3][0] ), .IN4(n144), .Q(
          n198));
   AO22X1 U194 (.IN1(n346), .IN2(mem_write_data[1]), .IN3(\memory[3][1] ), .IN4(n144), .Q(
          n199));
   AO22X1 U195 (.IN1(n346), .IN2(mem_write_data[2]), .IN3(\memory[3][2] ), .IN4(n144), .Q(
          n200));
   AO22X1 U196 (.IN1(n346), .IN2(mem_write_data[3]), .IN3(\memory[3][3] ), .IN4(n144), .Q(
          n201));
   AO22X1 U197 (.IN1(n346), .IN2(mem_write_data[4]), .IN3(\memory[3][4] ), .IN4(n144), .Q(
          n202));
   AO22X1 U198 (.IN1(n346), .IN2(mem_write_data[5]), .IN3(\memory[3][5] ), .IN4(n144), .Q(
          n203));
   AO22X1 U199 (.IN1(n346), .IN2(mem_write_data[6]), .IN3(\memory[3][6] ), .IN4(n144), .Q(
          n204));
   AO22X1 U200 (.IN1(n346), .IN2(mem_write_data[7]), .IN3(\memory[3][7] ), .IN4(n144), .Q(
          n205));
   AO22X1 U201 (.IN1(n346), .IN2(mem_write_data[8]), .IN3(\memory[3][8] ), .IN4(n144), .Q(
          n206));
   AO22X1 U202 (.IN1(n346), .IN2(mem_write_data[9]), .IN3(\memory[3][9] ), .IN4(n144), .Q(
          n207));
   AO22X1 U203 (.IN1(n346), .IN2(mem_write_data[10]), .IN3(\memory[3][10] ), .IN4(n144), .
          Q(n208));
   AO22X1 U204 (.IN1(n346), .IN2(mem_write_data[11]), .IN3(\memory[3][11] ), .IN4(n144), .
          Q(n209));
   AO22X1 U205 (.IN1(n346), .IN2(mem_write_data[12]), .IN3(\memory[3][12] ), .IN4(n144), .
          Q(n210));
   AO22X1 U206 (.IN1(n346), .IN2(mem_write_data[13]), .IN3(\memory[3][13] ), .IN4(n144), .
          Q(n211));
   AO22X1 U207 (.IN1(n346), .IN2(mem_write_data[14]), .IN3(\memory[3][14] ), .IN4(n144), .
          Q(n212));
   AO22X1 U208 (.IN1(n346), .IN2(mem_write_data[15]), .IN3(\memory[3][15] ), .IN4(n144), .
          Q(n213));
   AO22X1 U210 (.IN1(n353), .IN2(mem_write_data[0]), .IN3(\memory[4][0] ), .IN4(n145), .Q(
          n214));
   AO22X1 U211 (.IN1(n353), .IN2(mem_write_data[1]), .IN3(\memory[4][1] ), .IN4(n145), .Q(
          n215));
   AO22X1 U212 (.IN1(n353), .IN2(mem_write_data[2]), .IN3(\memory[4][2] ), .IN4(n145), .Q(
          n216));
   AO22X1 U213 (.IN1(n353), .IN2(mem_write_data[3]), .IN3(\memory[4][3] ), .IN4(n145), .Q(
          n217));
   AO22X1 U214 (.IN1(n353), .IN2(mem_write_data[4]), .IN3(\memory[4][4] ), .IN4(n145), .Q(
          n218));
   AO22X1 U215 (.IN1(n353), .IN2(mem_write_data[5]), .IN3(\memory[4][5] ), .IN4(n145), .Q(
          n219));
   AO22X1 U216 (.IN1(n353), .IN2(mem_write_data[6]), .IN3(\memory[4][6] ), .IN4(n145), .Q(
          n220));
   AO22X1 U217 (.IN1(n353), .IN2(mem_write_data[7]), .IN3(\memory[4][7] ), .IN4(n145), .Q(
          n221));
   AO22X1 U218 (.IN1(n353), .IN2(mem_write_data[8]), .IN3(\memory[4][8] ), .IN4(n145), .Q(
          n222));
   AO22X1 U219 (.IN1(n353), .IN2(mem_write_data[9]), .IN3(\memory[4][9] ), .IN4(n145), .Q(
          n223));
   AO22X1 U220 (.IN1(n353), .IN2(mem_write_data[10]), .IN3(\memory[4][10] ), .IN4(n145), .
          Q(n224));
   AO22X1 U221 (.IN1(n353), .IN2(mem_write_data[11]), .IN3(\memory[4][11] ), .IN4(n145), .
          Q(n225));
   AO22X1 U222 (.IN1(n353), .IN2(mem_write_data[12]), .IN3(\memory[4][12] ), .IN4(n145), .
          Q(n226));
   AO22X1 U223 (.IN1(n353), .IN2(mem_write_data[13]), .IN3(\memory[4][13] ), .IN4(n145), .
          Q(n227));
   AO22X1 U224 (.IN1(n353), .IN2(mem_write_data[14]), .IN3(\memory[4][14] ), .IN4(n145), .
          Q(n228));
   AO22X1 U225 (.IN1(n353), .IN2(mem_write_data[15]), .IN3(\memory[4][15] ), .IN4(n145), .
          Q(n229));
   AO22X1 U227 (.IN1(n352), .IN2(mem_write_data[0]), .IN3(\memory[5][0] ), .IN4(n147), .Q(
          n230));
   AO22X1 U228 (.IN1(n352), .IN2(mem_write_data[1]), .IN3(\memory[5][1] ), .IN4(n147), .Q(
          n231));
   AO22X1 U229 (.IN1(n352), .IN2(mem_write_data[2]), .IN3(\memory[5][2] ), .IN4(n147), .Q(
          n232));
   AO22X1 U230 (.IN1(n352), .IN2(mem_write_data[3]), .IN3(\memory[5][3] ), .IN4(n147), .Q(
          n233));
   AO22X1 U231 (.IN1(n352), .IN2(mem_write_data[4]), .IN3(\memory[5][4] ), .IN4(n147), .Q(
          n234));
   AO22X1 U232 (.IN1(n352), .IN2(mem_write_data[5]), .IN3(\memory[5][5] ), .IN4(n147), .Q(
          n235));
   AO22X1 U233 (.IN1(n352), .IN2(mem_write_data[6]), .IN3(\memory[5][6] ), .IN4(n147), .Q(
          n236));
   AO22X1 U234 (.IN1(n352), .IN2(mem_write_data[7]), .IN3(\memory[5][7] ), .IN4(n147), .Q(
          n237));
   AO22X1 U235 (.IN1(n352), .IN2(mem_write_data[8]), .IN3(\memory[5][8] ), .IN4(n147), .Q(
          n238));
   AO22X1 U236 (.IN1(n352), .IN2(mem_write_data[9]), .IN3(\memory[5][9] ), .IN4(n147), .Q(
          n239));
   AO22X1 U237 (.IN1(n352), .IN2(mem_write_data[10]), .IN3(\memory[5][10] ), .IN4(n147), .
          Q(n240));
   AO22X1 U238 (.IN1(n352), .IN2(mem_write_data[11]), .IN3(\memory[5][11] ), .IN4(n147), .
          Q(n241));
   AO22X1 U239 (.IN1(n352), .IN2(mem_write_data[12]), .IN3(\memory[5][12] ), .IN4(n147), .
          Q(n242));
   AO22X1 U240 (.IN1(n352), .IN2(mem_write_data[13]), .IN3(\memory[5][13] ), .IN4(n147), .
          Q(n243));
   AO22X1 U241 (.IN1(n352), .IN2(mem_write_data[14]), .IN3(\memory[5][14] ), .IN4(n147), .
          Q(n244));
   AO22X1 U242 (.IN1(n352), .IN2(mem_write_data[15]), .IN3(\memory[5][15] ), .IN4(n147), .
          Q(n245));
   AO22X1 U244 (.IN1(n351), .IN2(mem_write_data[0]), .IN3(\memory[6][0] ), .IN4(n148), .Q(
          n246));
   AO22X1 U245 (.IN1(n351), .IN2(mem_write_data[1]), .IN3(\memory[6][1] ), .IN4(n148), .Q(
          n247));
   AO22X1 U246 (.IN1(n351), .IN2(mem_write_data[2]), .IN3(\memory[6][2] ), .IN4(n148), .Q(
          n248));
   AO22X1 U247 (.IN1(n351), .IN2(mem_write_data[3]), .IN3(\memory[6][3] ), .IN4(n148), .Q(
          n249));
   AO22X1 U248 (.IN1(n351), .IN2(mem_write_data[4]), .IN3(\memory[6][4] ), .IN4(n148), .Q(
          n250));
   AO22X1 U249 (.IN1(n351), .IN2(mem_write_data[5]), .IN3(\memory[6][5] ), .IN4(n148), .Q(
          n251));
   AO22X1 U250 (.IN1(n351), .IN2(mem_write_data[6]), .IN3(\memory[6][6] ), .IN4(n148), .Q(
          n252));
   AO22X1 U251 (.IN1(n351), .IN2(mem_write_data[7]), .IN3(\memory[6][7] ), .IN4(n148), .Q(
          n253));
   AO22X1 U252 (.IN1(n351), .IN2(mem_write_data[8]), .IN3(\memory[6][8] ), .IN4(n148), .Q(
          n254));
   AO22X1 U253 (.IN1(n351), .IN2(mem_write_data[9]), .IN3(\memory[6][9] ), .IN4(n148), .Q(
          n255));
   AO22X1 U254 (.IN1(n351), .IN2(mem_write_data[10]), .IN3(\memory[6][10] ), .IN4(n148), .
          Q(n256));
   AO22X1 U255 (.IN1(n351), .IN2(mem_write_data[11]), .IN3(\memory[6][11] ), .IN4(n148), .
          Q(n257));
   AO22X1 U256 (.IN1(n351), .IN2(mem_write_data[12]), .IN3(\memory[6][12] ), .IN4(n148), .
          Q(n258));
   AO22X1 U257 (.IN1(n351), .IN2(mem_write_data[13]), .IN3(\memory[6][13] ), .IN4(n148), .
          Q(n259));
   AO22X1 U258 (.IN1(n351), .IN2(mem_write_data[14]), .IN3(\memory[6][14] ), .IN4(n148), .
          Q(n260));
   AO22X1 U259 (.IN1(n351), .IN2(mem_write_data[15]), .IN3(\memory[6][15] ), .IN4(n148), .
          Q(n261));
   AO22X1 U261 (.IN1(n350), .IN2(mem_write_data[0]), .IN3(\memory[7][0] ), .IN4(n344), .Q(
          n262));
   AO22X1 U262 (.IN1(n350), .IN2(mem_write_data[1]), .IN3(\memory[7][1] ), .IN4(n345), .Q(
          n263));
   AO22X1 U263 (.IN1(n350), .IN2(mem_write_data[2]), .IN3(\memory[7][2] ), .IN4(n344), .Q(
          n264));
   AO22X1 U264 (.IN1(n350), .IN2(mem_write_data[3]), .IN3(\memory[7][3] ), .IN4(n345), .Q(
          n265));
   AO22X1 U265 (.IN1(n350), .IN2(mem_write_data[4]), .IN3(\memory[7][4] ), .IN4(n344), .Q(
          n266));
   AO22X1 U266 (.IN1(n350), .IN2(mem_write_data[5]), .IN3(\memory[7][5] ), .IN4(n345), .Q(
          n267));
   AO22X1 U267 (.IN1(n350), .IN2(mem_write_data[6]), .IN3(\memory[7][6] ), .IN4(n344), .Q(
          n268));
   AO22X1 U268 (.IN1(n350), .IN2(mem_write_data[7]), .IN3(\memory[7][7] ), .IN4(n345), .Q(
          n269));
   AO22X1 U269 (.IN1(n350), .IN2(mem_write_data[8]), .IN3(\memory[7][8] ), .IN4(n344), .Q(
          n270));
   AO22X1 U270 (.IN1(n350), .IN2(mem_write_data[9]), .IN3(\memory[7][9] ), .IN4(n345), .Q(
          n271));
   AO22X1 U271 (.IN1(n350), .IN2(mem_write_data[10]), .IN3(\memory[7][10] ), .IN4(n344), .
          Q(n272));
   AO22X1 U272 (.IN1(n350), .IN2(mem_write_data[11]), .IN3(\memory[7][11] ), .IN4(n345), .
          Q(n273));
   AO22X1 U273 (.IN1(n350), .IN2(mem_write_data[12]), .IN3(\memory[7][12] ), .IN4(n344), .
          Q(n274));
   AO22X1 U274 (.IN1(n350), .IN2(mem_write_data[13]), .IN3(\memory[7][13] ), .IN4(n345), .
          Q(n275));
   AO22X1 U275 (.IN1(n350), .IN2(mem_write_data[14]), .IN3(\memory[7][14] ), .IN4(n344), .
          Q(n276));
   AO22X1 U276 (.IN1(n350), .IN2(mem_write_data[15]), .IN3(\memory[7][15] ), .IN4(n345), .
          Q(n277));
   AND2X1 U278 (.IN1(N14), .IN2(mem_write_en), .Q(n146));
   AND2X1 U279 (.IN1(mem_read), .IN2(N39), .Q(mem_read_data[9]));
   AND2X1 U280 (.IN1(N40), .IN2(mem_read), .Q(mem_read_data[8]));
   AND2X1 U281 (.IN1(N41), .IN2(mem_read), .Q(mem_read_data[7]));
   AND2X1 U282 (.IN1(N42), .IN2(mem_read), .Q(mem_read_data[6]));
   AND2X1 U283 (.IN1(N43), .IN2(mem_read), .Q(mem_read_data[5]));
   AND2X1 U284 (.IN1(N44), .IN2(mem_read), .Q(mem_read_data[4]));
   AND2X1 U285 (.IN1(N45), .IN2(mem_read), .Q(mem_read_data[3]));
   AND2X1 U286 (.IN1(N46), .IN2(mem_read), .Q(mem_read_data[2]));
   AND2X1 U287 (.IN1(N47), .IN2(mem_read), .Q(mem_read_data[1]));
   AND2X1 U288 (.IN1(N33), .IN2(mem_read), .Q(mem_read_data[15]));
   AND2X1 U289 (.IN1(N34), .IN2(mem_read), .Q(mem_read_data[14]));
   AND2X1 U290 (.IN1(N35), .IN2(mem_read), .Q(mem_read_data[13]));
   AND2X1 U291 (.IN1(N36), .IN2(mem_read), .Q(mem_read_data[12]));
   AND2X1 U292 (.IN1(N37), .IN2(mem_read), .Q(mem_read_data[11]));
   AND2X1 U293 (.IN1(N38), .IN2(mem_read), .Q(mem_read_data[10]));
   AND2X1 U294 (.IN1(N48), .IN2(mem_read), .Q(mem_read_data[0]));
   INVX0 U130 (.INP(n140), .ZN(n349));
   INVX0 U131 (.INP(n143), .ZN(n347));
   INVX0 U132 (.INP(n148), .ZN(n351));
   INVX0 U133 (.INP(n145), .ZN(n353));
   INVX0 U134 (.INP(N13), .ZN(n343));
   AND2X1 U135 (.IN1(n133), .IN2(n354), .Q(n331));
   AND2X1 U136 (.IN1(n131), .IN2(n354), .Q(n334));
   AND2X1 U137 (.IN1(n132), .IN2(n354), .Q(n332));
   AND2X1 U138 (.IN1(n130), .IN2(n354), .Q(n335));
   INVX0 U139 (.INP(n142), .ZN(n348));
   INVX0 U140 (.INP(n144), .ZN(n346));
   INVX0 U141 (.INP(n147), .ZN(n352));
   INVX0 U158 (.INP(n149), .ZN(n350));
   NAND3X0 U175 (.IN1(n354), .IN2(n343), .IN3(n146), .QN(n145));
   NAND3X0 U192 (.IN1(N13), .IN2(n354), .IN3(n146), .QN(n148));
   NAND3X0 U209 (.IN1(n354), .IN2(n343), .IN3(n141), .QN(n140));
   NAND3X0 U226 (.IN1(n141), .IN2(n354), .IN3(N13), .QN(n143));
   NBUFFX2 U243 (.INP(n149), .Z(n344));
   NBUFFX2 U260 (.INP(n149), .Z(n345));
   AND2X1 U277 (.IN1(n133), .IN2(N12), .Q(n336));
   AND2X1 U295 (.IN1(n131), .IN2(N12), .Q(n339));
   AND2X1 U296 (.IN1(N12), .IN2(n132), .Q(n337));
   AND2X1 U297 (.IN1(n130), .IN2(N12), .Q(n340));
   INVX0 U298 (.INP(N12), .ZN(n354));
   NAND3X0 U299 (.IN1(n141), .IN2(n343), .IN3(N12), .QN(n142));
   NAND3X0 U300 (.IN1(N12), .IN2(n141), .IN3(N13), .QN(n144));
   NAND3X0 U301 (.IN1(N12), .IN2(n343), .IN3(n146), .QN(n147));
   NAND3X0 U302 (.IN1(N13), .IN2(N12), .IN3(n146), .QN(n149));
   NOR2X0 U303 (.IN1(n355), .IN2(N14), .QN(n141));
   INVX0 U304 (.INP(mem_write_en), .ZN(n355));
   NOR2X0 U305 (.IN1(N13), .IN2(N14), .QN(n130));
   NOR2X0 U306 (.IN1(n343), .IN2(N14), .QN(n131));
   AND2X1 U307 (.IN1(N14), .IN2(N13), .Q(n132));
   AND2X1 U308 (.IN1(N14), .IN2(n343), .Q(n133));
   AO22X1 U309 (.IN1(\memory[6][0] ), .IN2(n332), .IN3(\memory[4][0] ), .IN4(n331), .Q(
          n129));
   AO221X1 U310 (.IN1(\memory[0][0] ), .IN2(n335), .IN3(\memory[2][0] ), .IN4(n334), .IN5(
          n129), .Q(n136));
   AO22X1 U311 (.IN1(\memory[7][0] ), .IN2(n337), .IN3(\memory[5][0] ), .IN4(n336), .Q(
          n134));
   AO221X1 U312 (.IN1(\memory[1][0] ), .IN2(n340), .IN3(\memory[3][0] ), .IN4(n339), .IN5(
          n134), .Q(n135));
   OR2X1 U313 (.IN1(n136), .IN2(n135), .Q(N48));
   AO22X1 U314 (.IN1(\memory[6][1] ), .IN2(n332), .IN3(\memory[4][1] ), .IN4(n331), .Q(
          n137));
   AO221X1 U315 (.IN1(\memory[0][1] ), .IN2(n335), .IN3(\memory[2][1] ), .IN4(n334), .IN5(
          n137), .Q(n278));
   AO22X1 U316 (.IN1(\memory[7][1] ), .IN2(n337), .IN3(\memory[5][1] ), .IN4(n336), .Q(
          n138));
   AO221X1 U317 (.IN1(\memory[1][1] ), .IN2(n340), .IN3(\memory[3][1] ), .IN4(n339), .IN5(
          n138), .Q(n139));
   OR2X1 U318 (.IN1(n278), .IN2(n139), .Q(N47));
   AO22X1 U319 (.IN1(\memory[6][2] ), .IN2(n332), .IN3(\memory[4][2] ), .IN4(n331), .Q(
          n279));
   AO221X1 U320 (.IN1(\memory[0][2] ), .IN2(n335), .IN3(\memory[2][2] ), .IN4(n334), .IN5(
          n279), .Q(n282));
   AO22X1 U321 (.IN1(\memory[7][2] ), .IN2(n337), .IN3(\memory[5][2] ), .IN4(n336), .Q(
          n280));
   AO221X1 U322 (.IN1(\memory[1][2] ), .IN2(n340), .IN3(\memory[3][2] ), .IN4(n339), .IN5(
          n280), .Q(n281));
   OR2X1 U323 (.IN1(n282), .IN2(n281), .Q(N46));
   AO22X1 U324 (.IN1(\memory[6][3] ), .IN2(n332), .IN3(\memory[4][3] ), .IN4(n331), .Q(
          n283));
   AO221X1 U325 (.IN1(\memory[0][3] ), .IN2(n335), .IN3(\memory[2][3] ), .IN4(n334), .IN5(
          n283), .Q(n286));
   AO22X1 U326 (.IN1(\memory[7][3] ), .IN2(n337), .IN3(\memory[5][3] ), .IN4(n336), .Q(
          n284));
   AO221X1 U327 (.IN1(\memory[1][3] ), .IN2(n340), .IN3(\memory[3][3] ), .IN4(n339), .IN5(
          n284), .Q(n285));
   OR2X1 U328 (.IN1(n286), .IN2(n285), .Q(N45));
   AO22X1 U329 (.IN1(\memory[6][4] ), .IN2(n332), .IN3(\memory[4][4] ), .IN4(n331), .Q(
          n287));
   AO221X1 U330 (.IN1(\memory[0][4] ), .IN2(n335), .IN3(\memory[2][4] ), .IN4(n334), .IN5(
          n287), .Q(n290));
   AO22X1 U331 (.IN1(\memory[7][4] ), .IN2(n337), .IN3(\memory[5][4] ), .IN4(n336), .Q(
          n288));
   AO221X1 U332 (.IN1(\memory[1][4] ), .IN2(n340), .IN3(\memory[3][4] ), .IN4(n339), .IN5(
          n288), .Q(n289));
   OR2X1 U333 (.IN1(n290), .IN2(n289), .Q(N44));
   AO22X1 U334 (.IN1(\memory[6][5] ), .IN2(n332), .IN3(\memory[4][5] ), .IN4(n331), .Q(
          n291));
   AO221X1 U335 (.IN1(\memory[0][5] ), .IN2(n335), .IN3(\memory[2][5] ), .IN4(n334), .IN5(
          n291), .Q(n294));
   AO22X1 U336 (.IN1(\memory[7][5] ), .IN2(n337), .IN3(\memory[5][5] ), .IN4(n336), .Q(
          n292));
   AO221X1 U337 (.IN1(\memory[1][5] ), .IN2(n340), .IN3(\memory[3][5] ), .IN4(n339), .IN5(
          n292), .Q(n293));
   OR2X1 U338 (.IN1(n294), .IN2(n293), .Q(N43));
   AO22X1 U339 (.IN1(\memory[6][6] ), .IN2(n332), .IN3(\memory[4][6] ), .IN4(n331), .Q(
          n295));
   AO221X1 U340 (.IN1(\memory[0][6] ), .IN2(n335), .IN3(\memory[2][6] ), .IN4(n334), .IN5(
          n295), .Q(n298));
   AO22X1 U341 (.IN1(\memory[7][6] ), .IN2(n337), .IN3(\memory[5][6] ), .IN4(n336), .Q(
          n296));
   AO221X1 U342 (.IN1(\memory[1][6] ), .IN2(n340), .IN3(\memory[3][6] ), .IN4(n339), .IN5(
          n296), .Q(n297));
   OR2X1 U343 (.IN1(n298), .IN2(n297), .Q(N42));
   AO22X1 U344 (.IN1(\memory[6][7] ), .IN2(n332), .IN3(\memory[4][7] ), .IN4(n331), .Q(
          n299));
   AO221X1 U345 (.IN1(\memory[0][7] ), .IN2(n335), .IN3(\memory[2][7] ), .IN4(n334), .IN5(
          n299), .Q(n302));
   AO22X1 U346 (.IN1(\memory[7][7] ), .IN2(n337), .IN3(\memory[5][7] ), .IN4(n336), .Q(
          n300));
   AO221X1 U347 (.IN1(\memory[1][7] ), .IN2(n340), .IN3(\memory[3][7] ), .IN4(n339), .IN5(
          n300), .Q(n301));
   OR2X1 U348 (.IN1(n302), .IN2(n301), .Q(N41));
   AO22X1 U349 (.IN1(\memory[6][8] ), .IN2(n332), .IN3(\memory[4][8] ), .IN4(n331), .Q(
          n303));
   AO221X1 U350 (.IN1(\memory[0][8] ), .IN2(n335), .IN3(\memory[2][8] ), .IN4(n334), .IN5(
          n303), .Q(n306));
   AO22X1 U351 (.IN1(\memory[7][8] ), .IN2(n337), .IN3(\memory[5][8] ), .IN4(n336), .Q(
          n304));
   AO221X1 U352 (.IN1(\memory[1][8] ), .IN2(n340), .IN3(\memory[3][8] ), .IN4(n339), .IN5(
          n304), .Q(n305));
   OR2X1 U353 (.IN1(n306), .IN2(n305), .Q(N40));
   AO22X1 U354 (.IN1(\memory[6][9] ), .IN2(n332), .IN3(\memory[4][9] ), .IN4(n331), .Q(
          n307));
   AO221X1 U355 (.IN1(\memory[0][9] ), .IN2(n335), .IN3(\memory[2][9] ), .IN4(n334), .IN5(
          n307), .Q(n310));
   AO22X1 U356 (.IN1(\memory[7][9] ), .IN2(n337), .IN3(\memory[5][9] ), .IN4(n336), .Q(
          n308));
   AO221X1 U357 (.IN1(\memory[1][9] ), .IN2(n340), .IN3(\memory[3][9] ), .IN4(n339), .IN5(
          n308), .Q(n309));
   OR2X1 U358 (.IN1(n310), .IN2(n309), .Q(N39));
   AO22X1 U359 (.IN1(\memory[6][10] ), .IN2(n332), .IN3(\memory[4][10] ), .IN4(n331), .Q(
          n311));
   AO221X1 U360 (.IN1(\memory[0][10] ), .IN2(n335), .IN3(\memory[2][10] ), .IN4(n334), .
          IN5(n311), .Q(n314));
   AO22X1 U361 (.IN1(\memory[7][10] ), .IN2(n337), .IN3(\memory[5][10] ), .IN4(n336), .Q(
          n312));
   AO221X1 U362 (.IN1(\memory[1][10] ), .IN2(n340), .IN3(\memory[3][10] ), .IN4(n339), .
          IN5(n312), .Q(n313));
   OR2X1 U363 (.IN1(n314), .IN2(n313), .Q(N38));
   AO22X1 U364 (.IN1(\memory[6][11] ), .IN2(n332), .IN3(\memory[4][11] ), .IN4(n331), .Q(
          n315));
   AO221X1 U365 (.IN1(\memory[0][11] ), .IN2(n335), .IN3(\memory[2][11] ), .IN4(n334), .
          IN5(n315), .Q(n318));
   AO22X1 U366 (.IN1(\memory[7][11] ), .IN2(n337), .IN3(\memory[5][11] ), .IN4(n336), .Q(
          n316));
   AO221X1 U367 (.IN1(\memory[1][11] ), .IN2(n340), .IN3(\memory[3][11] ), .IN4(n339), .
          IN5(n316), .Q(n317));
   OR2X1 U368 (.IN1(n318), .IN2(n317), .Q(N37));
   AO22X1 U369 (.IN1(\memory[6][12] ), .IN2(n332), .IN3(\memory[4][12] ), .IN4(n331), .Q(
          n319));
   AO221X1 U370 (.IN1(\memory[0][12] ), .IN2(n335), .IN3(\memory[2][12] ), .IN4(n334), .
          IN5(n319), .Q(n322));
   AO22X1 U371 (.IN1(\memory[7][12] ), .IN2(n337), .IN3(\memory[5][12] ), .IN4(n336), .Q(
          n320));
   AO221X1 U372 (.IN1(\memory[1][12] ), .IN2(n340), .IN3(\memory[3][12] ), .IN4(n339), .
          IN5(n320), .Q(n321));
   OR2X1 U373 (.IN1(n322), .IN2(n321), .Q(N36));
   AO22X1 U374 (.IN1(\memory[6][13] ), .IN2(n332), .IN3(\memory[4][13] ), .IN4(n331), .Q(
          n323));
   AO221X1 U375 (.IN1(\memory[0][13] ), .IN2(n335), .IN3(\memory[2][13] ), .IN4(n334), .
          IN5(n323), .Q(n326));
   AO22X1 U376 (.IN1(\memory[7][13] ), .IN2(n337), .IN3(\memory[5][13] ), .IN4(n336), .Q(
          n324));
   AO221X1 U377 (.IN1(\memory[1][13] ), .IN2(n340), .IN3(\memory[3][13] ), .IN4(n339), .
          IN5(n324), .Q(n325));
   OR2X1 U378 (.IN1(n326), .IN2(n325), .Q(N35));
   AO22X1 U379 (.IN1(\memory[6][14] ), .IN2(n332), .IN3(\memory[4][14] ), .IN4(n331), .Q(
          n327));
   AO221X1 U380 (.IN1(\memory[0][14] ), .IN2(n335), .IN3(\memory[2][14] ), .IN4(n334), .
          IN5(n327), .Q(n330));
   AO22X1 U381 (.IN1(\memory[7][14] ), .IN2(n337), .IN3(\memory[5][14] ), .IN4(n336), .Q(
          n328));
   AO221X1 U382 (.IN1(\memory[1][14] ), .IN2(n340), .IN3(\memory[3][14] ), .IN4(n339), .
          IN5(n328), .Q(n329));
   OR2X1 U383 (.IN1(n330), .IN2(n329), .Q(N34));
   AO22X1 U384 (.IN1(\memory[6][15] ), .IN2(n332), .IN3(\memory[4][15] ), .IN4(n331), .Q(
          n333));
   AO221X1 U385 (.IN1(\memory[0][15] ), .IN2(n335), .IN3(\memory[2][15] ), .IN4(n334), .
          IN5(n333), .Q(n342));
   AO22X1 U386 (.IN1(\memory[7][15] ), .IN2(n337), .IN3(\memory[5][15] ), .IN4(n336), .Q(
          n338));
   AO221X1 U387 (.IN1(\memory[1][15] ), .IN2(n340), .IN3(\memory[3][15] ), .IN4(n339), .
          IN5(n338), .Q(n341));
   OR2X1 U388 (.IN1(n342), .IN2(n341), .Q(N33));
endmodule

module Datapath_Unit_test_1 (clk, jump, beq, mem_read, mem_write, alu_src, reg_dst, 
       mem_to_reg, reg_write, bne, alu_op, opcode, test_si3, test_si2, test_si1, test_so3
       , test_so2, test_so1, test_se);
input clk, jump, beq, mem_read, mem_write, alu_src, reg_dst, mem_to_reg, reg_write, bne, 
       test_si3, test_si2, test_si1, test_se;
input [1:0] alu_op;
output test_so3, test_so2, test_so1;
output [3:0] opcode;
wire zero_flag, n28, n29, n30, \add_37/carry[15] , \add_37/carry[14] , \add_37/carry[13] 
       , \add_37/carry[12] , \add_37/carry[11] , \add_37/carry[10] , \add_37/carry[9] , 
       \add_37/carry[8] , \add_37/carry[7] , \add_37/carry[6] , \add_37/carry[5] , 
       \add_37/carry[4] , \add_37/carry[3] , n1, n2, n3, n4, n5, n22, n23, n24, n25, n26, 
       n27, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
       , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n63, 
       n64, n65, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83
       , n84;
wire [15:0] pc_current;
wire [15:0] pc_next;
wire [11:0] instr;
wire [15:0] reg_write_data;
wire [15:0] reg_read_data_1;
wire [15:0] reg_read_data_2;
wire [2:0] ALU_Control;
wire [15:0] ALU_out;
wire [15:0] PC_2beq;
wire [15:0] mem_read_data;
   assign opcode[3] = 1'b0;
   assign opcode[2] = 1'b0;
   assign opcode[1] = 1'b0;
   assign opcode[0] = 1'b0;
   SDFFX1 \pc_current_reg[0]  (.D(pc_next[0]), .SI(n84), .SE(test_se), .CLK(clk), .Q(
          PC_2beq[0]), .QN(n83));
   SDFFX1 \pc_current_reg[15]  (.D(pc_next[15]), .SI(n70), .SE(test_se), .CLK(clk), .Q(
          pc_current[15]), .QN(n69));
   SDFFX1 \pc_current_reg[9]  (.D(pc_next[9]), .SI(n76), .SE(test_se), .CLK(clk), .Q(
          pc_current[9]), .QN(n75));
   SDFFX1 \pc_current_reg[8]  (.D(pc_next[8]), .SI(n77), .SE(test_se), .CLK(clk), .Q(
          pc_current[8]), .QN(n76));
   SDFFX1 \pc_current_reg[7]  (.D(pc_next[7]), .SI(n78), .SE(test_se), .CLK(clk), .Q(
          pc_current[7]), .QN(n77));
   SDFFX1 \pc_current_reg[6]  (.D(pc_next[6]), .SI(n79), .SE(test_se), .CLK(clk), .Q(
          pc_current[6]), .QN(n78));
   SDFFX1 \pc_current_reg[5]  (.D(pc_next[5]), .SI(n80), .SE(test_se), .CLK(clk), .Q(
          pc_current[5]), .QN(n79));
   SDFFX1 \pc_current_reg[4]  (.D(pc_next[4]), .SI(n81), .SE(test_se), .CLK(clk), .Q(
          pc_current[4]), .QN(n80));
   SDFFX1 \pc_current_reg[3]  (.D(pc_next[3]), .SI(n82), .SE(test_se), .CLK(clk), .Q(
          pc_current[3]), .QN(n81));
   SDFFX1 \pc_current_reg[2]  (.D(pc_next[2]), .SI(n1), .SE(test_se), .CLK(clk), .Q(
          pc_current[2]), .QN(n82));
   SDFFX1 \pc_current_reg[1]  (.D(pc_next[1]), .SI(n83), .SE(test_se), .CLK(clk), .Q(
          pc_current[1]), .QN(n1));
   SDFFX1 \pc_current_reg[14]  (.D(pc_next[14]), .SI(n71), .SE(test_se), .CLK(clk), .Q(
          pc_current[14]), .QN(n70));
   SDFFX1 \pc_current_reg[13]  (.D(pc_next[13]), .SI(n72), .SE(test_se), .CLK(clk), .Q(
          pc_current[13]), .QN(n71));
   SDFFX1 \pc_current_reg[12]  (.D(pc_next[12]), .SI(n73), .SE(test_se), .CLK(clk), .Q(
          pc_current[12]), .QN(n72));
   SDFFX1 \pc_current_reg[11]  (.D(pc_next[11]), .SI(n74), .SE(test_se), .CLK(clk), .Q(
          pc_current[11]), .QN(n73));
   SDFFX1 \pc_current_reg[10]  (.D(pc_next[10]), .SI(n75), .SE(test_se), .CLK(clk), .Q(
          pc_current[10]), .QN(n74));
   AO22X1 U32 (.IN1(mem_to_reg), .IN2(mem_read_data[9]), .IN3(ALU_out[9]), .IN4(n37), .Q(
          reg_write_data[9]));
   AO22X1 U33 (.IN1(mem_read_data[8]), .IN2(mem_to_reg), .IN3(ALU_out[8]), .IN4(n37), .Q(
          reg_write_data[8]));
   AO22X1 U34 (.IN1(mem_read_data[7]), .IN2(mem_to_reg), .IN3(ALU_out[7]), .IN4(n37), .Q(
          reg_write_data[7]));
   AO22X1 U35 (.IN1(mem_read_data[6]), .IN2(mem_to_reg), .IN3(ALU_out[6]), .IN4(n37), .Q(
          reg_write_data[6]));
   AO22X1 U36 (.IN1(mem_read_data[5]), .IN2(mem_to_reg), .IN3(ALU_out[5]), .IN4(n37), .Q(
          reg_write_data[5]));
   AO22X1 U37 (.IN1(mem_read_data[4]), .IN2(mem_to_reg), .IN3(ALU_out[4]), .IN4(n37), .Q(
          reg_write_data[4]));
   AO22X1 U38 (.IN1(mem_read_data[3]), .IN2(mem_to_reg), .IN3(ALU_out[3]), .IN4(n37), .Q(
          reg_write_data[3]));
   AO22X1 U39 (.IN1(mem_read_data[2]), .IN2(mem_to_reg), .IN3(ALU_out[2]), .IN4(n37), .Q(
          reg_write_data[2]));
   AO22X1 U40 (.IN1(mem_read_data[1]), .IN2(mem_to_reg), .IN3(ALU_out[1]), .IN4(n37), .Q(
          reg_write_data[1]));
   AO22X1 U41 (.IN1(mem_read_data[15]), .IN2(mem_to_reg), .IN3(ALU_out[15]), .IN4(n37), .Q(
          reg_write_data[15]));
   AO22X1 U42 (.IN1(mem_read_data[14]), .IN2(mem_to_reg), .IN3(ALU_out[14]), .IN4(n37), .Q(
          reg_write_data[14]));
   AO22X1 U43 (.IN1(mem_read_data[13]), .IN2(mem_to_reg), .IN3(ALU_out[13]), .IN4(n37), .Q(
          reg_write_data[13]));
   AO22X1 U44 (.IN1(mem_read_data[12]), .IN2(mem_to_reg), .IN3(ALU_out[12]), .IN4(n37), .Q(
          reg_write_data[12]));
   AO22X1 U45 (.IN1(mem_read_data[11]), .IN2(mem_to_reg), .IN3(ALU_out[11]), .IN4(n37), .Q(
          reg_write_data[11]));
   AO22X1 U46 (.IN1(mem_read_data[10]), .IN2(mem_to_reg), .IN3(ALU_out[10]), .IN4(n37), .Q(
          reg_write_data[10]));
   AO22X1 U47 (.IN1(mem_read_data[0]), .IN2(mem_to_reg), .IN3(ALU_out[0]), .IN4(n37), .Q(
          reg_write_data[0]));
   AO222X1 U74 (.IN1(PC_2beq[15]), .IN2(n28), .IN3(PC_2beq[15]), .IN4(n29), .IN5(
          PC_2beq[15]), .IN6(jump), .Q(pc_next[15]));
   AO222X1 U75 (.IN1(PC_2beq[14]), .IN2(n28), .IN3(PC_2beq[14]), .IN4(n29), .IN5(
          PC_2beq[14]), .IN6(jump), .Q(pc_next[14]));
   AO222X1 U76 (.IN1(PC_2beq[13]), .IN2(n28), .IN3(PC_2beq[13]), .IN4(n29), .IN5(
          PC_2beq[13]), .IN6(jump), .Q(pc_next[13]));
   AO22X1 U80 (.IN1(PC_2beq[0]), .IN2(n28), .IN3(PC_2beq[0]), .IN4(n29), .Q(pc_next[0]));
   Instruction_Memory im (.pc({pc_current[15:1], PC_2beq[0]}));
   GPRs_test_1 reg_file (.clk(clk), .reg_write_en(reg_write), .reg_write_dest({1'b0, 1'b0
          , 1'b0}), .reg_write_data(reg_write_data), .reg_read_addr_1({1'b0, 1'b0, 1'b0})
          , .reg_read_data_1(reg_read_data_1), .reg_read_addr_2({1'b0, 1'b0, 1'b0}), .
          reg_read_data_2(reg_read_data_2), .test_si2(test_si3), .test_si1(n69), .test_so2(
          test_so3), .test_so1(test_so2), .test_se(test_se));
   alu_control ALU_Control_unit (.ALU_Control(ALU_Control), .ALUOp(alu_op), .Function({
          1'b0, 1'b0, 1'b0, 1'b0}));
   ALU alu_unit (.a(reg_read_data_1), .b({n31, n23, n32, n36, n26, n24, n33, n27, n35, n25
          , n34, n3, n2, n22, n5, n4}), .alu_control(ALU_Control), .result(ALU_out), .zero(
          zero_flag));
   Data_Memory_test_1 dm (.clk(clk), .mem_access_addr(ALU_out), .mem_write_data(
          reg_read_data_2), .mem_write_en(mem_write), .mem_read(mem_read), .mem_read_data(
          mem_read_data), .test_si2(test_si2), .test_si1(test_si1), .test_so2(n84), .
          test_so1(test_so1), .test_se(test_se));
   AND2X1 U6 (.IN1(reg_read_data_2[3]), .IN2(n65), .Q(n2));
   AND2X1 U7 (.IN1(reg_read_data_2[4]), .IN2(n65), .Q(n3));
   NOR2X0 U21 (.IN1(n30), .IN2(jump), .QN(n29));
   NOR2X0 U22 (.IN1(n63), .IN2(jump), .QN(n28));
   INVX0 U23 (.INP(n30), .ZN(n63));
   INVX0 U24 (.INP(alu_src), .ZN(n65));
   AND2X1 U25 (.IN1(reg_read_data_2[0]), .IN2(n65), .Q(n4));
   AND2X1 U26 (.IN1(reg_read_data_2[1]), .IN2(n65), .Q(n5));
   AND2X1 U27 (.IN1(reg_read_data_2[2]), .IN2(n65), .Q(n22));
   AND2X1 U28 (.IN1(reg_read_data_2[14]), .IN2(n65), .Q(n23));
   AND2X1 U29 (.IN1(reg_read_data_2[10]), .IN2(n65), .Q(n24));
   AND2X1 U30 (.IN1(reg_read_data_2[6]), .IN2(n65), .Q(n25));
   AND2X1 U31 (.IN1(reg_read_data_2[11]), .IN2(n65), .Q(n26));
   AND2X1 U48 (.IN1(reg_read_data_2[8]), .IN2(n65), .Q(n27));
   AND2X1 U49 (.IN1(reg_read_data_2[15]), .IN2(n65), .Q(n31));
   AND2X1 U50 (.IN1(reg_read_data_2[13]), .IN2(n65), .Q(n32));
   AND2X1 U51 (.IN1(reg_read_data_2[9]), .IN2(n65), .Q(n33));
   AND2X1 U52 (.IN1(reg_read_data_2[5]), .IN2(n65), .Q(n34));
   AND2X1 U53 (.IN1(reg_read_data_2[7]), .IN2(n65), .Q(n35));
   AND2X1 U54 (.IN1(reg_read_data_2[12]), .IN2(n65), .Q(n36));
   NOR2X0 U55 (.IN1(n64), .IN2(zero_flag), .QN(n30));
   INVX0 U56 (.INP(bne), .ZN(n64));
   INVX0 U57 (.INP(mem_to_reg), .ZN(n37));
   NAND2X1 U58 (.IN1(n38), .IN2(n39), .QN(pc_next[12]));
   NAND2X1 U59 (.IN1(PC_2beq[12]), .IN2(n28), .QN(n38));
   NAND2X1 U60 (.IN1(PC_2beq[12]), .IN2(n29), .QN(n39));
   NAND2X1 U61 (.IN1(n40), .IN2(n41), .QN(pc_next[11]));
   NAND2X1 U62 (.IN1(PC_2beq[11]), .IN2(n28), .QN(n40));
   NAND2X1 U63 (.IN1(PC_2beq[11]), .IN2(n29), .QN(n41));
   NAND2X1 U64 (.IN1(n42), .IN2(n43), .QN(pc_next[10]));
   NAND2X1 U65 (.IN1(PC_2beq[10]), .IN2(n28), .QN(n42));
   NAND2X1 U66 (.IN1(PC_2beq[10]), .IN2(n29), .QN(n43));
   NAND2X1 U67 (.IN1(n44), .IN2(n45), .QN(pc_next[9]));
   NAND2X1 U68 (.IN1(PC_2beq[9]), .IN2(n28), .QN(n44));
   NAND2X1 U69 (.IN1(PC_2beq[9]), .IN2(n29), .QN(n45));
   NAND2X1 U70 (.IN1(n46), .IN2(n47), .QN(pc_next[8]));
   NAND2X1 U71 (.IN1(PC_2beq[8]), .IN2(n28), .QN(n46));
   NAND2X1 U72 (.IN1(PC_2beq[8]), .IN2(n29), .QN(n47));
   NAND2X1 U73 (.IN1(n48), .IN2(n49), .QN(pc_next[7]));
   NAND2X1 U77 (.IN1(PC_2beq[7]), .IN2(n28), .QN(n48));
   NAND2X1 U78 (.IN1(PC_2beq[7]), .IN2(n29), .QN(n49));
   NAND2X1 U79 (.IN1(n50), .IN2(n51), .QN(pc_next[6]));
   NAND2X1 U81 (.IN1(PC_2beq[6]), .IN2(n28), .QN(n50));
   NAND2X1 U82 (.IN1(PC_2beq[6]), .IN2(n29), .QN(n51));
   NAND2X1 U83 (.IN1(n52), .IN2(n53), .QN(pc_next[5]));
   NAND2X1 U84 (.IN1(PC_2beq[5]), .IN2(n28), .QN(n52));
   NAND2X1 U85 (.IN1(PC_2beq[5]), .IN2(n29), .QN(n53));
   NAND2X1 U86 (.IN1(n54), .IN2(n55), .QN(pc_next[4]));
   NAND2X1 U87 (.IN1(PC_2beq[4]), .IN2(n28), .QN(n54));
   NAND2X1 U88 (.IN1(PC_2beq[4]), .IN2(n29), .QN(n55));
   NAND2X1 U89 (.IN1(n56), .IN2(n57), .QN(pc_next[3]));
   NAND2X1 U90 (.IN1(PC_2beq[3]), .IN2(n28), .QN(n56));
   NAND2X1 U91 (.IN1(PC_2beq[3]), .IN2(n29), .QN(n57));
   NAND2X1 U92 (.IN1(n58), .IN2(n59), .QN(pc_next[2]));
   NAND2X1 U93 (.IN1(PC_2beq[2]), .IN2(n28), .QN(n58));
   NAND2X1 U94 (.IN1(PC_2beq[2]), .IN2(n29), .QN(n59));
   NAND2X1 U95 (.IN1(n60), .IN2(n61), .QN(pc_next[1]));
   NAND2X1 U96 (.IN1(n1), .IN2(n28), .QN(n60));
   NAND2X1 U97 (.IN1(n1), .IN2(n29), .QN(n61));
   XOR2X1 U98 (.IN1(pc_current[15]), .IN2(\add_37/carry[15] ), .Q(PC_2beq[15]));
   AND2X1 U99 (.IN1(pc_current[14]), .IN2(\add_37/carry[14] ), .Q(\add_37/carry[15] ));
   XOR2X1 U100 (.IN1(pc_current[14]), .IN2(\add_37/carry[14] ), .Q(PC_2beq[14]));
   AND2X1 U101 (.IN1(pc_current[13]), .IN2(\add_37/carry[13] ), .Q(\add_37/carry[14] ));
   XOR2X1 U102 (.IN1(pc_current[13]), .IN2(\add_37/carry[13] ), .Q(PC_2beq[13]));
   AND2X1 U103 (.IN1(pc_current[12]), .IN2(\add_37/carry[12] ), .Q(\add_37/carry[13] ));
   XOR2X1 U104 (.IN1(pc_current[12]), .IN2(\add_37/carry[12] ), .Q(PC_2beq[12]));
   AND2X1 U105 (.IN1(pc_current[11]), .IN2(\add_37/carry[11] ), .Q(\add_37/carry[12] ));
   XOR2X1 U106 (.IN1(pc_current[11]), .IN2(\add_37/carry[11] ), .Q(PC_2beq[11]));
   AND2X1 U107 (.IN1(pc_current[10]), .IN2(\add_37/carry[10] ), .Q(\add_37/carry[11] ));
   XOR2X1 U108 (.IN1(pc_current[10]), .IN2(\add_37/carry[10] ), .Q(PC_2beq[10]));
   AND2X1 U109 (.IN1(pc_current[9]), .IN2(\add_37/carry[9] ), .Q(\add_37/carry[10] ));
   XOR2X1 U110 (.IN1(pc_current[9]), .IN2(\add_37/carry[9] ), .Q(PC_2beq[9]));
   AND2X1 U111 (.IN1(pc_current[8]), .IN2(\add_37/carry[8] ), .Q(\add_37/carry[9] ));
   XOR2X1 U112 (.IN1(pc_current[8]), .IN2(\add_37/carry[8] ), .Q(PC_2beq[8]));
   AND2X1 U113 (.IN1(pc_current[7]), .IN2(\add_37/carry[7] ), .Q(\add_37/carry[8] ));
   XOR2X1 U114 (.IN1(pc_current[7]), .IN2(\add_37/carry[7] ), .Q(PC_2beq[7]));
   AND2X1 U115 (.IN1(pc_current[6]), .IN2(\add_37/carry[6] ), .Q(\add_37/carry[7] ));
   XOR2X1 U116 (.IN1(pc_current[6]), .IN2(\add_37/carry[6] ), .Q(PC_2beq[6]));
   AND2X1 U117 (.IN1(pc_current[5]), .IN2(\add_37/carry[5] ), .Q(\add_37/carry[6] ));
   XOR2X1 U118 (.IN1(pc_current[5]), .IN2(\add_37/carry[5] ), .Q(PC_2beq[5]));
   AND2X1 U119 (.IN1(pc_current[4]), .IN2(\add_37/carry[4] ), .Q(\add_37/carry[5] ));
   XOR2X1 U120 (.IN1(pc_current[4]), .IN2(\add_37/carry[4] ), .Q(PC_2beq[4]));
   AND2X1 U121 (.IN1(pc_current[3]), .IN2(\add_37/carry[3] ), .Q(\add_37/carry[4] ));
   XOR2X1 U122 (.IN1(pc_current[3]), .IN2(\add_37/carry[3] ), .Q(PC_2beq[3]));
   AND2X1 U123 (.IN1(pc_current[2]), .IN2(pc_current[1]), .Q(\add_37/carry[3] ));
   XOR2X1 U124 (.IN1(pc_current[2]), .IN2(pc_current[1]), .Q(PC_2beq[2]));
endmodule

module Control_Unit (opcode, alu_op, jump, beq, bne, mem_read, mem_write, alu_src, reg_dst
       , mem_to_reg, reg_write);
input [3:0] opcode;
output jump, beq, bne, mem_read, mem_write, alu_src, reg_dst, mem_to_reg, reg_write;
output [1:0] alu_op;
wire \alu_op[1] , n5, n6, n7, n8, n1, n2, n3, n4;
   assign alu_src = \alu_op[1] ;
   assign alu_op[1] = \alu_op[1] ;
   assign mem_to_reg = mem_read;
   AO21X1 U12 (.IN1(n1), .IN2(n4), .IN3(n5), .Q(reg_write));
   AO21X1 U13 (.IN1(opcode[1]), .IN2(n1), .IN3(n5), .Q(reg_dst));
   AO21X1 U14 (.IN1(opcode[2]), .IN2(opcode[1]), .IN3(n6), .Q(n5));
   XNOR2X1 U15 (.IN1(opcode[3]), .IN2(n7), .Q(n6));
   NOR3X0 U16 (.IN1(opcode[2]), .IN2(opcode[3]), .IN3(opcode[1]), .QN(\alu_op[1] ));
   OR2X1 U17 (.IN1(bne), .IN2(beq), .Q(alu_op[0]));
   AND4X1 U18 (.IN1(opcode[0]), .IN2(opcode[3]), .IN3(opcode[1]), .IN4(n4), .Q(beq));
   NAND3X0 U19 (.IN1(opcode[2]), .IN2(n2), .IN3(opcode[3]), .QN(n8));
   NOR2X0 U3 (.IN1(n1), .IN2(n8), .QN(jump));
   INVX0 U4 (.INP(\alu_op[1] ), .ZN(n3));
   NOR2X0 U5 (.IN1(n3), .IN2(n1), .QN(mem_write));
   NOR2X0 U6 (.IN1(opcode[0]), .IN2(n3), .QN(mem_read));
   NOR2X0 U7 (.IN1(n8), .IN2(opcode[0]), .QN(bne));
   NOR2X0 U8 (.IN1(opcode[1]), .IN2(opcode[2]), .QN(n7));
   INVX0 U9 (.INP(opcode[0]), .ZN(n1));
   INVX0 U10 (.INP(opcode[1]), .ZN(n2));
   INVX0 U11 (.INP(opcode[2]), .ZN(n4));
endmodule

module Risc_16_bit_DW01_add_width3 (A, B, CI, SUM, CO);
input CI;
input [2:0] A;
input [2:0] B;
output CO;
output [2:0] SUM;
wire n4, n5;
   NAND2X2 U1 (.IN1(B[0]), .IN2(A[0]), .QN(n5));
   XNOR2X1 U2 (.IN1(n4), .IN2(A[2]), .Q(SUM[2]));
   NAND3X0 U3 (.IN1(A[1]), .IN2(A[0]), .IN3(B[0]), .QN(n4));
   XNOR2X1 U4 (.IN1(A[1]), .IN2(n5), .Q(SUM[1]));
   XOR2X1 U5 (.IN1(B[0]), .IN2(A[0]), .Q(SUM[0]));
endmodule

module Risc_16_bit_DFT_cntr_scnto_width3_count_to5_rst_mode0_dcod_mode0_0_0
       (clk, rst_n, enable, load_n, tercnt_n, count);
input clk, rst_n, enable, load_n;
output tercnt_n;
output [2:0] count;
wire n6, n10, n9, n8, n13, n11, n14, n1;
   Risc_16_bit_DW01_add_width3 add_124 (.A(count), .B({1'b0, 1'b0, enable}), .CI(1'b0), .
          SUM({n10, n9, n8}));
   DFFARX1 \count_int_reg[0]  (.D(n11), .CLK(clk), .RSTB(rst_n), .Q(count[0]));
   DFFARX1 \count_int_reg[1]  (.D(n14), .CLK(clk), .RSTB(rst_n), .Q(count[1]));
   DFFARX1 \count_int_reg[2]  (.D(n13), .CLK(clk), .RSTB(rst_n), .Q(count[2]));
   DFFARX1 tercnt_n_reg_reg (.D(n6), .CLK(clk), .RSTB(rst_n), .QN(tercnt_n));
   INVX1 U4 (.INP(n9), .ZN(n1));
   AND3X1 U5 (.IN1(n8), .IN2(n1), .IN3(n13), .Q(n6));
   AND2X1 U6 (.IN1(load_n), .IN2(n9), .Q(n14));
   AND2X1 U7 (.IN1(n10), .IN2(load_n), .Q(n13));
   AND2X1 U8 (.IN1(load_n), .IN2(n8), .Q(n11));
endmodule

module Risc_16_bit_DFT_decode_width4_0_0 (A, B);
input [2:0] A;
output [7:0] B;
wire n1, n2, n3;
   INVX1 U2 (.INP(A[2]), .ZN(n1));
   INVX1 U3 (.INP(A[1]), .ZN(n2));
   INVX1 U4 (.INP(A[0]), .ZN(n3));
   AND3X1 U5 (.IN1(A[1]), .IN2(A[0]), .IN3(A[2]), .Q(B[7]));
   NOR3X0 U6 (.IN1(n1), .IN2(A[0]), .IN3(n2), .QN(B[6]));
   NOR3X0 U7 (.IN1(n1), .IN2(A[1]), .IN3(n3), .QN(B[5]));
   NOR3X0 U8 (.IN1(n1), .IN2(A[1]), .IN3(A[0]), .QN(B[4]));
   NOR3X0 U9 (.IN1(n2), .IN2(A[2]), .IN3(n3), .QN(B[3]));
   NOR3X0 U10 (.IN1(n2), .IN2(A[2]), .IN3(A[0]), .QN(B[2]));
   NOR3X0 U11 (.IN1(n3), .IN2(A[2]), .IN3(A[1]), .QN(B[1]));
   NOR3X0 U12 (.IN1(A[0]), .IN2(A[2]), .IN3(A[1]), .QN(B[0]));
endmodule

module Risc_16_bit_DFT_or_gate_width4_0_0 (a, b);
input [3:0] a;
output b;
   OR4X1 U1 (.IN1(a[1]), .IN2(a[0]), .IN3(a[3]), .IN4(a[2]), .Q(b));
endmodule

module Risc_16_bit_DFT_clk_control_0_0 (reset, scan_en, clk_enable, fast_clk, slow_clk, 
       fast_clk_enable, slow_clk_enable);
input reset, scan_en, fast_clk, slow_clk;
input [3:0] clk_enable;
output fast_clk_enable, slow_clk_enable;
wire n5, n6, n10, n9, n8, n7, n15, n14, n13, n12, n21, n20, n19, n22, n23, n25, n26, n28, 
       n29, n31, n1, n2, n3, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
       SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
   Risc_16_bit_DFT_cntr_scnto_width3_count_to5_rst_mode0_dcod_mode0_0_0 U_cycle_ctr_i
          (.clk(fast_clk), .rst_n(n2), .enable(n22), .load_n(n25), .tercnt_n(n23), .count({
          n21, n20, n19}));
   Risc_16_bit_DFT_decode_width4_0_0 U_decode_i (.A({n21, n20, n19}), .B({
          SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, n15, 
          n14, n13, n12, SYNOPSYS_UNCONNECTED__3}));
   Risc_16_bit_DFT_or_gate_width4_0_0 U_or_tree_i (.a({n10, n9, n8, n7}), .b(n6));
   DFFARX1 pipeline_or_tree_l_reg (.D(n6), .CLK(fast_clk), .RSTB(n2), .Q(n5));
   DFFNARX1 fast_clk_enable_l_reg (.D(n31), .CLK(fast_clk), .RSTB(n2), .Q(fast_clk_enable)
          );
   DFFNARX1 slow_clk_enable_l_reg (.D(n29), .CLK(slow_clk), .RSTB(n2), .Q(slow_clk_enable)
          , .QN(n1));
   DFFARX1 load_n_meta_0_l_reg (.D(n1), .CLK(fast_clk), .RSTB(n2), .Q(n28));
   DFFARX1 load_n_meta_1_l_reg (.D(n28), .CLK(fast_clk), .RSTB(n2), .Q(n26));
   DFFARX1 load_n_meta_2_l_reg (.D(n26), .CLK(fast_clk), .RSTB(n2), .Q(n25));
   NOR2X2 U3 (.IN1(fast_clk_enable), .IN2(n3), .QN(n29));
   INVX1 U4 (.INP(reset), .ZN(n2));
   INVX1 U5 (.INP(scan_en), .ZN(n3));
   AND2X1 U6 (.IN1(n14), .IN2(clk_enable[2]), .Q(n9));
   AND2X1 U7 (.IN1(n13), .IN2(clk_enable[1]), .Q(n8));
   AND2X1 U8 (.IN1(n12), .IN2(clk_enable[0]), .Q(n7));
   AND3X1 U9 (.IN1(n3), .IN2(n1), .IN3(n5), .Q(n31));
   AND2X1 U10 (.IN1(n23), .IN2(n3), .Q(n22));
   AND2X1 U11 (.IN1(n15), .IN2(clk_enable[3]), .Q(n10));
endmodule

module Risc_16_bit_DFT_gf_mux_0_0 (fast_clk_enable, slow_clk_enable, pll_bypass, test_mode
       , scan_en, fast_gate, slow_gate);
input fast_clk_enable, slow_clk_enable, pll_bypass, test_mode, scan_en;
output fast_gate, slow_gate;
wire n1, n2;
   OA21X2 U1 (.IN1(n2), .IN2(pll_bypass), .IN3(test_mode), .Q(slow_gate));
   INVX1 U2 (.INP(fast_clk_enable), .ZN(n1));
   AND2X1 U3 (.IN1(slow_clk_enable), .IN2(scan_en), .Q(n2));
   OAI21X1 U4 (.IN1(n1), .IN2(pll_bypass), .IN3(test_mode), .QN(fast_gate));
endmodule

module Risc_16_bit_mselector_n2_m1_0 (DATA1_0, DATA2_0, CONTROL1, CONTROL2, Z_0);
input DATA1_0, DATA2_0, CONTROL1, CONTROL2;
output Z_0;
   AO22X1 U2 (.IN1(DATA2_0), .IN2(CONTROL2), .IN3(DATA1_0), .IN4(CONTROL1), .Q(Z_0));
endmodule

module Risc_16_bit_mselector_n2_m1 (DATA1_0, DATA2_0, CONTROL1, CONTROL2, Z_0);
input DATA1_0, DATA2_0, CONTROL1, CONTROL2;
output Z_0;
   AO22X1 U2 (.IN1(DATA2_0), .IN2(CONTROL2), .IN3(DATA1_0), .IN4(CONTROL1), .Q(Z_0));
endmodule

module Risc_16_bit_DFT_clk_mux_0 (fast_clk, scan_en, test_mode, reset, pll_bypass, 
       slow_clk, clk_enable, clk);
input fast_clk, scan_en, test_mode, reset, pll_bypass, slow_clk;
input [3:0] clk_enable;
output clk;
wire n6, n7, n21, n23, n2, n3, n4;
   Risc_16_bit_DFT_clk_control_0_0 U_clk_control_i_0 (.reset(reset), .scan_en(scan_en), .
          clk_enable(clk_enable), .fast_clk(fast_clk), .slow_clk(slow_clk), .
          fast_clk_enable(n7), .slow_clk_enable(n6));
   Risc_16_bit_DFT_gf_mux_0_0 U_gf_mux_0 (.fast_clk_enable(n7), .slow_clk_enable(n6), .
          pll_bypass(pll_bypass), .test_mode(test_mode), .scan_en(scan_en), .fast_gate(n23)
          , .slow_gate(n21));
   Risc_16_bit_mselector_n2_m1_0 U2 (.DATA1_0(fast_clk), .DATA2_0(n2), .CONTROL1(n23), .
          CONTROL2(n4), .Z_0(clk));
   Risc_16_bit_mselector_n2_m1 U3 (.DATA1_0(slow_clk), .DATA2_0(1'b0), .CONTROL1(n21), .
          CONTROL2(n3), .Z_0(n2));
   INVX1 U5 (.INP(n21), .ZN(n3));
   INVX1 U6 (.INP(n23), .ZN(n4));
endmodule

module Risc_16_bit_DFT_clk_chain_0 (clk, se, si, so, clk_ctrl_data);
input clk, se, si;
output so;
output [3:0] clk_ctrl_data;
wire n7, n14, n21, n28, n1;
   assign clk_ctrl_data[3] = so;
   DFFNX1 \U_shftreg_0/ff_3/q_reg  (.D(n28), .CLK(clk), .Q(clk_ctrl_data[0]));
   DFFNX1 \U_shftreg_0/ff_2/q_reg  (.D(n21), .CLK(clk), .Q(clk_ctrl_data[1]));
   DFFNX1 \U_shftreg_0/ff_1/q_reg  (.D(n14), .CLK(clk), .Q(clk_ctrl_data[2]));
   DFFNX1 \U_shftreg_0/ff_0/q_reg  (.D(n7), .CLK(clk), .Q(so));
   INVX1 U1 (.INP(se), .ZN(n1));
   AO22X1 U2 (.IN1(so), .IN2(n1), .IN3(se), .IN4(clk_ctrl_data[2]), .Q(n7));
   AO22X1 U3 (.IN1(si), .IN2(se), .IN3(clk_ctrl_data[0]), .IN4(n1), .Q(n28));
   AO22X1 U4 (.IN1(clk_ctrl_data[0]), .IN2(se), .IN3(clk_ctrl_data[1]), .IN4(n1), .Q(n21)
          );
   AO22X1 U5 (.IN1(clk_ctrl_data[2]), .IN2(n1), .IN3(clk_ctrl_data[1]), .IN4(se), .Q(n14)
          );
endmodule

module Risc_16_bit (clk, TEST_SI1, TEST_SI2, TEST_SI3, TEST_SI4, TEST_SE, TEST_SO1, 
       TEST_SO2, TEST_SO3, TEST_SO4, scan_clk, SCAN_MODE, pll_bypass_2, pll_bypass, 
       pll_reset);
input clk, TEST_SI1, TEST_SI2, TEST_SI3, TEST_SI4, TEST_SE, scan_clk, SCAN_MODE, 
       pll_bypass_2, pll_bypass, pll_reset;
output TEST_SO1, TEST_SO2, TEST_SO3, TEST_SO4;
wire n15, jump, beq, mem_read, mem_write, alu_src, reg_dst, mem_to_reg, reg_write, bne, n2
       , \clk_ctrl_data[0] , \clk_ctrl_data[1] , \clk_ctrl_data[2] , \clk_ctrl_data[3] , 
       n13;
wire [1:0] alu_op;
   Datapath_Unit_test_1 DU (.clk(n15), .jump(jump), .beq(beq), .mem_read(mem_read), .
          mem_write(mem_write), .alu_src(alu_src), .reg_dst(reg_dst), .mem_to_reg(n2), .
          reg_write(reg_write), .bne(bne), .alu_op(alu_op), .test_si3(TEST_SI4), .test_si2(
          TEST_SI3), .test_si1(TEST_SI1), .test_so3(TEST_SO4), .test_so2(TEST_SO3), .
          test_so1(TEST_SO1), .test_se(TEST_SE));
   Control_Unit control (.opcode({1'b0, 1'b0, 1'b0, 1'b0}), .alu_op(alu_op), .jump(jump), .
          beq(beq), .bne(bne), .mem_read(mem_read), .mem_write(mem_write), .alu_src(
          alu_src), .reg_dst(reg_dst), .mem_to_reg(mem_to_reg), .reg_write(reg_write));
   NBUFFX2 U1 (.INP(mem_to_reg), .Z(n2));
   Risc_16_bit_DFT_clk_mux_0 occ_snps_pll_controller (.fast_clk(clk), .scan_en(TEST_SE), .
          test_mode(n13), .reset(pll_reset), .pll_bypass(pll_bypass), .slow_clk(scan_clk)
          , .clk_enable({\clk_ctrl_data[3] , \clk_ctrl_data[2] , \clk_ctrl_data[1] , 
          \clk_ctrl_data[0] }), .clk(n15));
   Risc_16_bit_DFT_clk_chain_0 snps_clk_chain_0 (.clk(n15), .se(TEST_SE), .si(TEST_SI2), .
          so(TEST_SO2), .clk_ctrl_data({\clk_ctrl_data[3] , \clk_ctrl_data[2] , 
          \clk_ctrl_data[1] , \clk_ctrl_data[0] }));
   INVX0 U3 (.INP(SCAN_MODE), .ZN(n13));
endmodule

