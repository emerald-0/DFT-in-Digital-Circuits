// Verilog netlist written by  TetraMAX(R)  U-2022.12-SP7-i20231010_191200 
// Date: Mon May 20 15:22:02 2024

module LSDNENX1 (ENB, D, Q);
input ENB, D;
output Q;
   or or0 (Q, ENB, D);
endmodule

module SDFFSSRX2 (CLK, D, RSTB, SETB, SI, SE, Q, QN);
input CLK, D, RSTB, SETB, SI, SE;
output Q, QN;
wire S, DS, D1, D2, Q_buf, setb, rstb, nD, nCLK, nSE, nSI, CLK_D_RSTB_SI_SE, RSTB_CLK_D, 
       CLK_nD_RSTB_nSI_nSE, RSTB_nCLK_D, RSTB_nCLK_nD, CLK_D_SETB_SI_SE, 
       CLK_nD_SETB_nSI_nSE, nCLK_D_SETB, nCLK_nD_SETB, D_RSTB_SI_SE, nD_RSTB_nSI_nSE, 
       CLK_D_RSTB, RSTB_CLK_nD, nCLK_D_RSTB, nCLK_nD_RSTB, D_SETB, nD_SETB, CLK_D_SETB, 
       CLK_nD_SETB, CLK_D, CLK_RSTB, CLK_SETB, CLK_nD, nCLK_D, nCLK_nD, D_SE, D_SI, D_RSTB
       , RSTB_SETB, RSTB_D_SETB, RSTB_nD_SETB, RSTB_nD, RSTB_i, SETB_i, CLK_check, D_check
       ;
reg notifier;
   pullup pullup0 (setb);
   pullup pullup1 (rstb);
   not not2 (S, SETB);
   or or3 (DS, S, D);
   and and4 (D1, DS, RSTB);
   saed90_mux saed90_mux5 (D2, D1, SI, SE);
   saed90_dff_pos saed90_dff_pos6 (Q_buf, D2, CLK, rstb, setb, notifier);
   buf buf7 (Q, Q_buf);
   not not8 (QN, Q_buf);
   not not9 (nD, D);
   not not10 (nCLK, CLK);
   not not11 (nSE, SE);
   not not12 (nSI, SI);
   and and13 (CLK_D_RSTB_SI_SE, CLK, D, RSTB, SI, SE);
   and and14 (RSTB_CLK_D, RSTB, CLK, D);
   and and15 (CLK_nD_RSTB_nSI_nSE, CLK, nD, RSTB, nSI, nSE);
   and and16 (RSTB_nCLK_D, RSTB, nCLK, D);
   and and17 (RSTB_nCLK_nD, RSTB, nCLK, nD);
   and and18 (CLK_D_SETB_SI_SE, CLK, D, SETB, SI, SE);
   and and19 (CLK_nD_SETB_nSI_nSE, CLK, nD, SETB, nSI, nSE);
   and and20 (nCLK_D_SETB, nCLK, D, SETB);
   and and21 (nCLK_nD_SETB, nCLK, nD, SETB);
   and and22 (D_RSTB_SI_SE, D, RSTB, SI, SE);
   and and23 (nD_RSTB_nSI_nSE, nD, RSTB, nSI, nSE);
   and and24 (CLK_D_RSTB, CLK, D, RSTB);
   and and25 (RSTB_CLK_nD, RSTB, CLK, nD);
   and and26 (nCLK_D_RSTB, nCLK, D, RSTB);
   and and27 (nCLK_nD_RSTB, nCLK, nD, RSTB);
   and and28 (D_SETB, D, SETB);
   and and29 (nD_SETB, nD, SETB);
   and and30 (CLK_D_SETB, CLK, D, SETB);
   and and31 (CLK_nD_SETB, CLK, nD, SETB);
   and and32 (nCLK_D_SETB, nCLK, D, SETB);
   and and33 (nCLK_nD_SETB, nCLK, nD, SETB);
   and and34 (CLK_D, CLK, D);
   and and35 (CLK_RSTB, CLK, RSTB);
   and and36 (CLK_SETB, CLK, SETB);
   and and37 (CLK_nD, CLK, nD);
   and and38 (nCLK_D, nCLK, D);
   and and39 (nCLK_nD, nCLK, nD);
   and and40 (D_SE, D, SE);
   and and41 (D_SI, D, SI);
   and and42 (D_RSTB, D, RSTB);
   and and43 (D_SETB, D, SETB);
   and and44 (RSTB_SETB, RSTB, SETB);
   and and45 (RSTB_D_SETB, RSTB, D, SETB);
   and and46 (RSTB_nD_SETB, RSTB, nD, SETB);
   and and47 (RSTB_nD, RSTB, nD);
   buf buf48 (RSTB_i, RSTB);
   buf buf49 (SETB_i, SETB);
   and and50 (CLK_check, RSTB_i, SETB_i);
   and and51 (D_check, RSTB_i, SETB_i);
endmodule

`suppress_faults
`enable_portfaults
module TIEL (ZN);
output ZN;
   buf buf0 (ZN, 1'b0);
endmodule
`disable_portfaults
`nosuppress_faults

module aes_encipher_block_test_1 (clk, reset_n, next, keylen, round, round_key, sboxw, 
       new_sboxw, block, new_block, ready, test_si, test_so, test_se);
input clk, reset_n, next, keylen, test_si, test_se;
input [127:0] round_key;
input [31:0] new_sboxw;
input [127:0] block;
output ready, test_so;
output [3:0] round;
output [31:0] sboxw;
output [127:0] new_block;
wire n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
       n171, n172, n173, n174, n175, n177, n178, n179, n180, n181, n182, n183, n184, n185
       , n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
       n199, n200, n201, n202, n203, n204, n206, n207, n208, n209, n210, n211, n213, n214
       , n215, n216, n217, n218, n219, n220, n221, n223, n224, n225, n226, n227, n228, 
       n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n275
       , n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
       n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302
       , n303, n304, n305, n306, n307, n308, n309, n310, n312, n313, n314, n315, n316, 
       n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330
       , n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
       n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357
       , n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
       n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n384, n385
       , n386, n387, n388, n389, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
       n400, n401, n402, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414
       , n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
       n428, n429, n430, n431, n432, n434, n435, n436, n437, n438, n439, n441, n442, n443
       , n444, n445, n446, n447, n448, n449, n450, n451, n452, n454, n455, n456, n457, 
       n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471
       , n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n484, n485, 
       n486, n487, n488, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500
       , n502, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, 
       n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529
       , n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
       n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556
       , n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
       n570, n571, n573, n574, n575, n576, n577, n578, n580, n581, n582, n583, n584, n585
       , n586, n587, n588, n589, n590, n591, n593, n594, n595, n596, n597, n598, n599, 
       n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613
       , n614, n615, n616, n617, n618, n619, n620, n621, n623, n624, n625, n626, n627, 
       n628, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n643
       , n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, 
       n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670
       , n671, n673, n674, n675, n676, n677, n679, n680, n681, n682, n683, n684, n685, 
       n686, n687, n688, n689, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700
       , n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
       n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728
       , n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
       n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755
       , n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, 
       n769, n771, n772, n773, n774, n775, n776, n778, n779, n780, n781, n782, n783, n784
       , n785, n786, n787, n788, n789, n791, n792, n793, n794, n795, n796, n797, n798, 
       n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812
       , n813, n814, n815, n816, n817, n818, n819, n821, n822, n823, n824, n825, n826, 
       n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n841, n842
       , n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
       n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869
       , n871, n872, n873, n874, n875, n877, n878, n879, n880, n881, n882, n883, n884, 
       n885, n886, n887, n889, n890, n891, n892, n893, n894, n895, n896, n898, n899, n900
       , n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, 
       n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927
       , n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, 
       n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954
       , n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n967, n968, 
       n969, n970, n971, n972, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983
       , n984, n985, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, 
       n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
       n1010, n1011, n1012, n1013, n1014, n1015, n1017, n1018, n1019, n1020, n1021, n1022
       , n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, 
       n1035, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047
       , n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
       n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1067, n1068, n1069, n1070, n1071
       , n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
       n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096
       , n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
       n1108, n1109, n1110, n1111, n1112, n1114, n1115, n1116, n1117, n1118, n1119, n1120
       , n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
       n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143
       , n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
       n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166
       , n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, 
       n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189
       , n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, 
       n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212
       , n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
       n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235
       , n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
       n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1, n2, n3, n4, n142, n143, n144, 
       n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n176, n205
       , n212, n222, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
       n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266
       , n267, n268, n269, n270, n271, n272, n273, n274, n311, n383, n390, n403, n433, 
       n440, n453, n483, n489, n501, n503, n572, n579, n592, n622, n629, n642, n672, n678
       , n690, n701, n770, n777, n790, n820, n827, n840, n870, n876, n888, n897, n966, 
       n973, n986, n1016, n1023, n1036, n1066, n1072, n1084, n1113, n1254, n1255, n1256, 
       n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268
       , n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
       n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291
       , n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
       n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314
       , n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1323, n1324, n1325, n1326, 
       n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338
       , n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
       n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361
       , n1362;
wire [1:0] sword_ctr_reg;
wire [1:0] enc_ctrl_reg;
   assign test_so = n179;
   SDFFARX1 \sword_ctr_reg_reg[0]  (.D(n1253), .SI(n175), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(sword_ctr_reg[0]), .QN(n180));
   SDFFARX1 \sword_ctr_reg_reg[1]  (.D(n1252), .SI(n180), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(sword_ctr_reg[1]), .QN(n179));
   SDFFARX1 \round_ctr_reg_reg[0]  (.D(n1249), .SI(n1323), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(round[0]), .QN(n178));
   SDFFARX1 \round_ctr_reg_reg[1]  (.D(n1248), .SI(n178), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(round[1]), .QN(n177));
   SDFFARX1 \round_ctr_reg_reg[2]  (.D(n1247), .SI(n177), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(round[2]), .QN(n274));
   SDFFARX1 \round_ctr_reg_reg[3]  (.D(n1246), .SI(n274), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(round[3]), .QN(n175));
   SDFFARX1 \enc_ctrl_reg_reg[1]  (.D(n1251), .SI(n158), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(enc_ctrl_reg[1]), .QN(n157));
   SDFFASX1 ready_reg_reg (.D(n1245), .SI(enc_ctrl_reg[1]), .SE(test_se), .CLK(clk), .SETB(
          n1278), .Q(ready), .QN(n1323));
   SDFFARX1 \block_w0_reg_reg[0]  (.D(n1244), .SI(test_si), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(new_block[96]), .QN(n1362));
   SDFFARX1 \block_w1_reg_reg[24]  (.D(n1155), .SI(n273), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(new_block[88]), .QN(n1341));
   SDFFARX1 \block_w1_reg_reg[16]  (.D(n1163), .SI(n1349), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(new_block[80]), .QN(n1348));
   SDFFARX1 \block_w0_reg_reg[17]  (.D(n1131), .SI(n1361), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(new_block[113]), .QN(n227));
   SDFFARX1 \block_w3_reg_reg[26]  (.D(n1217), .SI(n250), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[26]), .QN(n1327));
   SDFFARX1 \block_w3_reg_reg[18]  (.D(n1225), .SI(n165), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[18]), .QN(n164));
   SDFFARX1 \block_w2_reg_reg[26]  (.D(n1185), .SI(n260), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[58]), .QN(n184));
   SDFFARX1 \block_w2_reg_reg[18]  (.D(n1193), .SI(n191), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[50]), .QN(n190));
   SDFFARX1 \block_w1_reg_reg[26]  (.D(n1153), .SI(n252), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[90]), .QN(n1340));
   SDFFARX1 \block_w1_reg_reg[18]  (.D(n1161), .SI(n1347), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[82]), .QN(n1346));
   SDFFARX1 \block_w0_reg_reg[26]  (.D(n1122), .SI(n221), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[122]), .QN(n220));
   SDFFARX1 \block_w0_reg_reg[18]  (.D(n1130), .SI(n227), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[114]), .QN(n1360));
   SDFFARX1 \block_w3_reg_reg[19]  (.D(n1224), .SI(n164), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[19]), .QN(n163));
   SDFFARX1 \block_w2_reg_reg[11]  (.D(n1200), .SI(n194), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[43]), .QN(n193));
   SDFFARX1 \block_w0_reg_reg[12]  (.D(n1136), .SI(n232), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[108]), .QN(n231));
   SDFFARX1 \block_w2_reg_reg[28]  (.D(n1183), .SI(n258), .SE(test_se), .CLK(clk), .RSTB(
          n1268), .Q(new_block[60]), .QN(n151));
   SDFFARX1 \block_w2_reg_reg[29]  (.D(n1182), .SI(n151), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[61]), .QN(n183));
   SDFFARX1 \block_w2_reg_reg[21]  (.D(n1190), .SI(n188), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[53]), .QN(n187));
   SDFFARX1 \block_w1_reg_reg[30]  (.D(n1149), .SI(n206), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[94]), .QN(n1339));
   SDFFARX1 \block_w1_reg_reg[7]  (.D(n1172), .SI(n1353), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[71]), .QN(n269));
   SDFFARX1 \block_w2_reg_reg[31]  (.D(n1180), .SI(n182), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[63]), .QN(n181));
   SDFFARX1 \block_w2_reg_reg[24]  (.D(n1187), .SI(n185), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[56]), .QN(n1335));
   SDFFARX1 \block_w2_reg_reg[16]  (.D(n1195), .SI(n192), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[48]), .QN(n1336));
   SDFFARX1 \block_w1_reg_reg[17]  (.D(n1162), .SI(n1348), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[81]), .QN(n1347));
   SDFFARX1 \block_w0_reg_reg[25]  (.D(n1123), .SI(n1358), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[121]), .QN(n221));
   SDFFARX1 \block_w0_reg_reg[9]  (.D(n1139), .SI(n235), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[105]), .QN(n234));
   SDFFARX1 \block_w2_reg_reg[25]  (.D(n1186), .SI(n1335), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[57]), .QN(n260));
   SDFFARX1 \block_w2_reg_reg[17]  (.D(n1194), .SI(n1336), .SE(test_se), .CLK(clk), .RSTB(
          n1269), .Q(new_block[49]), .QN(n191));
   SDFFARX1 \block_w1_reg_reg[25]  (.D(n1154), .SI(n1341), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[89]), .QN(n252));
   SDFFARX1 \block_w1_reg_reg[9]  (.D(n1170), .SI(n211), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[73]), .QN(n210));
   SDFFARX1 \block_w3_reg_reg[25]  (.D(n1218), .SI(n1328), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[25]), .QN(n250));
   SDFFARX1 \block_w3_reg_reg[17]  (.D(n1226), .SI(n1329), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[17]), .QN(n165));
   SDFFARX1 \block_w2_reg_reg[9]  (.D(n1202), .SI(n196), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[41]), .QN(n195));
   SDFFARX1 \block_w0_reg_reg[10]  (.D(n1138), .SI(n234), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[106]), .QN(n233));
   SDFFARX1 \block_w2_reg_reg[19]  (.D(n1192), .SI(n190), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[51]), .QN(n189));
   SDFFARX1 \block_w1_reg_reg[11]  (.D(n1168), .SI(n1352), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[75]), .QN(n209));
   SDFFARX1 \block_w3_reg_reg[12]  (.D(n1231), .SI(n167), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[12]), .QN(n176));
   SDFFARX1 \block_w1_reg_reg[28]  (.D(n1151), .SI(n256), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[92]), .QN(n207));
   SDFFARX1 \block_w1_reg_reg[5]  (.D(n1174), .SI(n214), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[69]), .QN(n213));
   SDFFARX1 \block_w2_reg_reg[14]  (.D(n1197), .SI(n1338), .SE(test_se), .CLK(clk), .RSTB(
          n1270), .Q(new_block[46]), .QN(n1337));
   SDFFARX1 \block_w0_reg_reg[30]  (.D(n1118), .SI(n219), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[126]), .QN(n218));
   SDFFARX1 \block_w0_reg_reg[31]  (.D(n1117), .SI(n218), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[127]), .QN(n1355));
   SDFFARX1 \block_w0_reg_reg[24]  (.D(n1124), .SI(n1359), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[120]), .QN(n1358));
   SDFFARX1 \block_w0_reg_reg[16]  (.D(n1132), .SI(n228), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[112]), .QN(n1361));
   SDFFARX1 \block_w3_reg_reg[24]  (.D(n1219), .SI(n159), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[24]), .QN(n1328));
   SDFFARX1 \block_w3_reg_reg[16]  (.D(n1227), .SI(n166), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[16]), .QN(n1329));
   SDFFARX1 \block_w2_reg_reg[8]  (.D(n1203), .SI(n197), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[40]), .QN(n196));
   SDFFARX1 \block_w0_reg_reg[8]  (.D(n1140), .SI(n236), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[104]), .QN(n235));
   SDFFARX1 \block_w2_reg_reg[0]  (.D(n1211), .SI(n268), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[32]), .QN(n204));
   SDFFARX1 \block_w3_reg_reg[1]  (.D(n1242), .SI(n1334), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[1]), .QN(n271));
   SDFFARX1 \block_w0_reg_reg[2]  (.D(n1146), .SI(n262), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[98]), .QN(n241));
   SDFFARX1 \block_w1_reg_reg[10]  (.D(n1169), .SI(n210), .SE(test_se), .CLK(clk), .RSTB(
          n1271), .Q(new_block[74]), .QN(n1352));
   SDFFARX1 \block_w3_reg_reg[11]  (.D(n1232), .SI(n168), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[11]), .QN(n167));
   SDFFARX1 \block_w1_reg_reg[27]  (.D(n1152), .SI(n1340), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[91]), .QN(n256));
   SDFFARX1 \block_w1_reg_reg[19]  (.D(n1160), .SI(n1346), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[83]), .QN(n1345));
   SDFFARX1 \block_w0_reg_reg[27]  (.D(n1121), .SI(n220), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[123]), .QN(n1357));
   SDFFARX1 \block_w0_reg_reg[19]  (.D(n1129), .SI(n1360), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[115]), .QN(n226));
   SDFFARX1 \block_w3_reg_reg[27]  (.D(n1216), .SI(n1327), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[27]), .QN(n244));
   SDFFARX1 \block_w3_reg_reg[4]  (.D(n1239), .SI(n173), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[4]), .QN(n172));
   SDFFARX1 \block_w0_reg_reg[28]  (.D(n1120), .SI(n1357), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[124]), .QN(n1356));
   SDFFARX1 \block_w0_reg_reg[29]  (.D(n1119), .SI(n1356), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[125]), .QN(n219));
   SDFFARX1 \block_w0_reg_reg[21]  (.D(n1127), .SI(n225), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[117]), .QN(n224));
   SDFFARX1 \block_w3_reg_reg[30]  (.D(n1213), .SI(n1326), .SE(test_se), .CLK(clk), .RSTB(
          n1272), .Q(new_block[30]), .QN(n1325));
   SDFFARX1 \block_w3_reg_reg[31]  (.D(n1212), .SI(n1325), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[31]), .QN(n1324));
   SDFFARX1 \block_w3_reg_reg[23]  (.D(n1220), .SI(n160), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[23]), .QN(n159));
   SDFFARX1 \block_w2_reg_reg[23]  (.D(n1188), .SI(n186), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[55]), .QN(n185));
   SDFFARX1 \block_w1_reg_reg[15]  (.D(n1164), .SI(n1350), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[79]), .QN(n1349));
   SDFFARX1 \block_w3_reg_reg[15]  (.D(n1228), .SI(n1330), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[15]), .QN(n166));
   SDFFARX1 \block_w1_reg_reg[12]  (.D(n1167), .SI(n209), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[76]), .QN(n208));
   SDFFARX1 \block_w3_reg_reg[21]  (.D(n1222), .SI(n162), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[21]), .QN(n161));
   SDFFARX1 \block_w2_reg_reg[30]  (.D(n1181), .SI(n183), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[62]), .QN(n182));
   SDFFARX1 \block_w2_reg_reg[22]  (.D(n1189), .SI(n187), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[54]), .QN(n186));
   SDFFARX1 \block_w1_reg_reg[31]  (.D(n1148), .SI(n1339), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[95]), .QN(n268));
   SDFFARX1 \block_w1_reg_reg[23]  (.D(n1156), .SI(n1342), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[87]), .QN(n273));
   SDFFARX1 \block_w0_reg_reg[23]  (.D(n1125), .SI(n223), .SE(test_se), .CLK(clk), .RSTB(
          n1273), .Q(new_block[119]), .QN(n1359));
   SDFFARX1 \block_w3_reg_reg[20]  (.D(n1223), .SI(n163), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[20]), .QN(n162));
   SDFFARX1 \block_w2_reg_reg[12]  (.D(n1199), .SI(n193), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[44]), .QN(n265));
   SDFFARX1 \block_w0_reg_reg[20]  (.D(n1128), .SI(n226), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[116]), .QN(n225));
   SDFFARX1 \block_w3_reg_reg[29]  (.D(n1214), .SI(n147), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[29]), .QN(n1326));
   SDFFARX1 \block_w3_reg_reg[13]  (.D(n1230), .SI(n176), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[13]), .QN(n1331));
   SDFFARX1 \block_w1_reg_reg[29]  (.D(n1150), .SI(n207), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[93]), .QN(n206));
   SDFFARX1 \block_w1_reg_reg[6]  (.D(n1173), .SI(n213), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[70]), .QN(n1353));
   SDFFARX1 \block_w2_reg_reg[15]  (.D(n1196), .SI(n1337), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[47]), .QN(n192));
   SDFFARX1 \block_w0_reg_reg[11]  (.D(n1137), .SI(n233), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[107]), .QN(n232));
   SDFFARX1 \block_w2_reg_reg[27]  (.D(n1184), .SI(n184), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[59]), .QN(n258));
   SDFFARX1 \block_w2_reg_reg[4]  (.D(n1207), .SI(n201), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[36]), .QN(n200));
   SDFFARX1 \block_w3_reg_reg[28]  (.D(n1215), .SI(n244), .SE(test_se), .CLK(clk), .RSTB(
          n1274), .Q(new_block[28]), .QN(n147));
   SDFFARX1 \block_w3_reg_reg[5]  (.D(n1238), .SI(n172), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[5]), .QN(n171));
   SDFFARX1 \block_w0_reg_reg[13]  (.D(n1135), .SI(n231), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[109]), .QN(n230));
   SDFFARX1 \block_w2_reg_reg[5]  (.D(n1206), .SI(n200), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[37]), .QN(n199));
   SDFFARX1 \block_w3_reg_reg[6]  (.D(n1237), .SI(n171), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[6]), .QN(n170));
   SDFFARX1 \block_w0_reg_reg[22]  (.D(n1126), .SI(n224), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[118]), .QN(n223));
   SDFFARX1 \block_w3_reg_reg[14]  (.D(n1229), .SI(n1331), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[14]), .QN(n1330));
   SDFFARX1 \block_w1_reg_reg[22]  (.D(n1157), .SI(n1343), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[86]), .QN(n1342));
   SDFFARX1 \block_w0_reg_reg[6]  (.D(n1142), .SI(n238), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[102]), .QN(n237));
   SDFFARX1 \block_w0_reg_reg[14]  (.D(n1134), .SI(n230), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[110]), .QN(n229));
   SDFFARX1 \block_w2_reg_reg[6]  (.D(n1205), .SI(n199), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[38]), .QN(n198));
   SDFFARX1 \block_w3_reg_reg[7]  (.D(n1236), .SI(n170), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[7]), .QN(n169));
   SDFFARX1 \block_w0_reg_reg[7]  (.D(n1141), .SI(n237), .SE(test_se), .CLK(clk), .RSTB(
          n1275), .Q(new_block[103]), .QN(n236));
   SDFFARX1 \block_w1_reg_reg[8]  (.D(n1171), .SI(n269), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[72]), .QN(n211));
   SDFFARX1 \block_w3_reg_reg[8]  (.D(n1235), .SI(n169), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[8]), .QN(n1333));
   SDFFARX1 \block_w1_reg_reg[0]  (.D(n1179), .SI(n1355), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[64]), .QN(n1354));
   SDFFARX1 \block_w0_reg_reg[15]  (.D(n1133), .SI(n229), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[111]), .QN(n228));
   SDFFARX1 \block_w2_reg_reg[7]  (.D(n1204), .SI(n198), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[39]), .QN(n197));
   SDFFARX1 \block_w3_reg_reg[0]  (.D(n1243), .SI(n181), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[0]), .QN(n1334));
   SDFFARX1 \block_w0_reg_reg[1]  (.D(n1147), .SI(n1362), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[97]), .QN(n262));
   SDFFARX1 \block_w1_reg_reg[1]  (.D(n1178), .SI(n1354), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[65]), .QN(n217));
   SDFFARX1 \block_w2_reg_reg[1]  (.D(n1210), .SI(n204), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[33]), .QN(n203));
   SDFFARX1 \block_w3_reg_reg[9]  (.D(n1234), .SI(n1333), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[9]), .QN(n1332));
   SDFFARX1 \block_w1_reg_reg[2]  (.D(n1177), .SI(n217), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[66]), .QN(n216));
   SDFFARX1 \block_w2_reg_reg[2]  (.D(n1209), .SI(n203), .SE(test_se), .CLK(clk), .RSTB(
          n1276), .Q(new_block[34]), .QN(n202));
   SDFFARX1 \block_w3_reg_reg[2]  (.D(n1241), .SI(n271), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[2]), .QN(n174));
   SDFFARX1 \block_w3_reg_reg[10]  (.D(n1233), .SI(n1332), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[10]), .QN(n168));
   SDFFARX1 \block_w2_reg_reg[10]  (.D(n1201), .SI(n195), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[42]), .QN(n194));
   SDFFARX1 \block_w2_reg_reg[3]  (.D(n1208), .SI(n202), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[35]), .QN(n201));
   SDFFARX1 \block_w3_reg_reg[3]  (.D(n1240), .SI(n174), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[3]), .QN(n173));
   SDFFARX1 \block_w0_reg_reg[3]  (.D(n1145), .SI(n241), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[99]), .QN(n240));
   SDFFARX1 \block_w1_reg_reg[3]  (.D(n1176), .SI(n216), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[67]), .QN(n215));
   SDFFARX1 \block_w2_reg_reg[20]  (.D(n1191), .SI(n189), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[52]), .QN(n188));
   SDFFARX1 \block_w1_reg_reg[20]  (.D(n1159), .SI(n1345), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[84]), .QN(n1344));
   SDFFARX1 \block_w0_reg_reg[4]  (.D(n1144), .SI(n240), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[100]), .QN(n239));
   SDFFARX1 \block_w1_reg_reg[4]  (.D(n1175), .SI(n215), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[68]), .QN(n214));
   SDFFARX1 \block_w2_reg_reg[13]  (.D(n1198), .SI(n265), .SE(test_se), .CLK(clk), .RSTB(
          n1277), .Q(new_block[45]), .QN(n1338));
   SDFFARX1 \block_w1_reg_reg[21]  (.D(n1158), .SI(n1344), .SE(test_se), .CLK(clk), .RSTB(
          n1278), .Q(new_block[85]), .QN(n1343));
   SDFFARX1 \block_w0_reg_reg[5]  (.D(n1143), .SI(n239), .SE(test_se), .CLK(clk), .RSTB(
          n1278), .Q(new_block[101]), .QN(n238));
   SDFFARX1 \block_w1_reg_reg[13]  (.D(n1166), .SI(n208), .SE(test_se), .CLK(clk), .RSTB(
          n1278), .Q(new_block[77]), .QN(n1351));
   SDFFARX1 \block_w1_reg_reg[14]  (.D(n1165), .SI(n1351), .SE(test_se), .CLK(clk), .RSTB(
          n1278), .Q(new_block[78]), .QN(n1350));
   SDFFARX1 \block_w3_reg_reg[22]  (.D(n1221), .SI(n161), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(new_block[22]), .QN(n160));
   AO221X1 U213 (.IN1(new_block[9]), .IN2(n489), .IN3(new_block[41]), .IN4(n383), .IN5(
          n275), .Q(sboxw[9]));
   AO22X1 U214 (.IN1(new_block[105]), .IN2(n572), .IN3(new_block[73]), .IN4(n440), .Q(n275)
          );
   AO221X1 U215 (.IN1(new_block[8]), .IN2(n1316), .IN3(new_block[40]), .IN4(n383), .IN5(
          n276), .Q(sboxw[8]));
   AO22X1 U216 (.IN1(new_block[104]), .IN2(n572), .IN3(new_block[72]), .IN4(n1315), .Q(
          n276));
   AO221X1 U217 (.IN1(new_block[7]), .IN2(n489), .IN3(new_block[39]), .IN4(n383), .IN5(
          n277), .Q(sboxw[7]));
   AO22X1 U218 (.IN1(new_block[103]), .IN2(n572), .IN3(new_block[71]), .IN4(n440), .Q(n277)
          );
   AO221X1 U219 (.IN1(new_block[6]), .IN2(n489), .IN3(new_block[38]), .IN4(n383), .IN5(
          n278), .Q(sboxw[6]));
   AO22X1 U220 (.IN1(new_block[102]), .IN2(n572), .IN3(new_block[70]), .IN4(n440), .Q(n278)
          );
   AO221X1 U221 (.IN1(new_block[5]), .IN2(n1316), .IN3(new_block[37]), .IN4(n383), .IN5(
          n279), .Q(sboxw[5]));
   AO22X1 U222 (.IN1(new_block[101]), .IN2(n572), .IN3(new_block[69]), .IN4(n1315), .Q(
          n279));
   AO221X1 U223 (.IN1(new_block[4]), .IN2(n489), .IN3(new_block[36]), .IN4(n383), .IN5(
          n280), .Q(sboxw[4]));
   AO22X1 U224 (.IN1(new_block[100]), .IN2(n572), .IN3(new_block[68]), .IN4(n440), .Q(n280)
          );
   AO221X1 U225 (.IN1(new_block[3]), .IN2(n489), .IN3(new_block[35]), .IN4(n383), .IN5(
          n281), .Q(sboxw[3]));
   AO22X1 U226 (.IN1(new_block[99]), .IN2(n572), .IN3(new_block[67]), .IN4(n440), .Q(n281)
          );
   AO221X1 U227 (.IN1(new_block[31]), .IN2(n489), .IN3(new_block[63]), .IN4(n383), .IN5(
          n282), .Q(sboxw[31]));
   AO22X1 U228 (.IN1(new_block[127]), .IN2(n572), .IN3(new_block[95]), .IN4(n440), .Q(n282)
          );
   AO221X1 U229 (.IN1(new_block[30]), .IN2(n489), .IN3(new_block[62]), .IN4(n383), .IN5(
          n283), .Q(sboxw[30]));
   AO22X1 U230 (.IN1(new_block[126]), .IN2(n572), .IN3(new_block[94]), .IN4(n440), .Q(n283)
          );
   AO221X1 U231 (.IN1(new_block[2]), .IN2(n489), .IN3(new_block[34]), .IN4(n383), .IN5(
          n284), .Q(sboxw[2]));
   AO22X1 U232 (.IN1(new_block[98]), .IN2(n572), .IN3(new_block[66]), .IN4(n440), .Q(n284)
          );
   AO221X1 U233 (.IN1(new_block[29]), .IN2(n1316), .IN3(new_block[61]), .IN4(n383), .IN5(
          n285), .Q(sboxw[29]));
   AO22X1 U234 (.IN1(new_block[125]), .IN2(n572), .IN3(new_block[93]), .IN4(n1315), .Q(
          n285));
   AO221X1 U235 (.IN1(new_block[28]), .IN2(n489), .IN3(new_block[60]), .IN4(n383), .IN5(
          n286), .Q(sboxw[28]));
   AO22X1 U236 (.IN1(new_block[124]), .IN2(n572), .IN3(new_block[92]), .IN4(n440), .Q(n286)
          );
   AO221X1 U237 (.IN1(new_block[27]), .IN2(n489), .IN3(new_block[59]), .IN4(n383), .IN5(
          n287), .Q(sboxw[27]));
   AO22X1 U238 (.IN1(new_block[123]), .IN2(n572), .IN3(new_block[91]), .IN4(n440), .Q(n287)
          );
   AO221X1 U239 (.IN1(new_block[26]), .IN2(n489), .IN3(new_block[58]), .IN4(n383), .IN5(
          n288), .Q(sboxw[26]));
   AO22X1 U240 (.IN1(new_block[122]), .IN2(n572), .IN3(new_block[90]), .IN4(n440), .Q(n288)
          );
   AO221X1 U241 (.IN1(new_block[25]), .IN2(n489), .IN3(new_block[57]), .IN4(n383), .IN5(
          n289), .Q(sboxw[25]));
   AO22X1 U242 (.IN1(new_block[121]), .IN2(n572), .IN3(new_block[89]), .IN4(n440), .Q(n289)
          );
   AO221X1 U243 (.IN1(new_block[24]), .IN2(n1316), .IN3(new_block[56]), .IN4(n383), .IN5(
          n290), .Q(sboxw[24]));
   AO22X1 U244 (.IN1(new_block[120]), .IN2(n572), .IN3(new_block[88]), .IN4(n1315), .Q(
          n290));
   AO221X1 U245 (.IN1(new_block[23]), .IN2(n489), .IN3(new_block[55]), .IN4(n383), .IN5(
          n291), .Q(sboxw[23]));
   AO22X1 U246 (.IN1(new_block[119]), .IN2(n572), .IN3(new_block[87]), .IN4(n440), .Q(n291)
          );
   AO221X1 U247 (.IN1(new_block[22]), .IN2(n489), .IN3(new_block[54]), .IN4(n383), .IN5(
          n292), .Q(sboxw[22]));
   AO22X1 U248 (.IN1(new_block[118]), .IN2(n572), .IN3(new_block[86]), .IN4(n440), .Q(n292)
          );
   AO221X1 U249 (.IN1(new_block[21]), .IN2(n1316), .IN3(new_block[53]), .IN4(n383), .IN5(
          n293), .Q(sboxw[21]));
   AO22X1 U250 (.IN1(new_block[117]), .IN2(n572), .IN3(new_block[85]), .IN4(n1315), .Q(
          n293));
   AO221X1 U251 (.IN1(new_block[20]), .IN2(n489), .IN3(new_block[52]), .IN4(n383), .IN5(
          n294), .Q(sboxw[20]));
   AO22X1 U252 (.IN1(new_block[116]), .IN2(n572), .IN3(new_block[84]), .IN4(n440), .Q(n294)
          );
   AO221X1 U253 (.IN1(new_block[1]), .IN2(n489), .IN3(new_block[33]), .IN4(n383), .IN5(
          n295), .Q(sboxw[1]));
   AO22X1 U254 (.IN1(new_block[97]), .IN2(n572), .IN3(new_block[65]), .IN4(n440), .Q(n295)
          );
   AO221X1 U255 (.IN1(new_block[19]), .IN2(n489), .IN3(new_block[51]), .IN4(n383), .IN5(
          n296), .Q(sboxw[19]));
   AO22X1 U256 (.IN1(new_block[115]), .IN2(n572), .IN3(new_block[83]), .IN4(n1315), .Q(
          n296));
   AO221X1 U257 (.IN1(new_block[18]), .IN2(n489), .IN3(new_block[50]), .IN4(n383), .IN5(
          n297), .Q(sboxw[18]));
   AO22X1 U258 (.IN1(new_block[114]), .IN2(n572), .IN3(new_block[82]), .IN4(n440), .Q(n297)
          );
   AO221X1 U259 (.IN1(new_block[17]), .IN2(n489), .IN3(new_block[49]), .IN4(n383), .IN5(
          n298), .Q(sboxw[17]));
   AO22X1 U260 (.IN1(new_block[113]), .IN2(n572), .IN3(new_block[81]), .IN4(n440), .Q(n298)
          );
   AO221X1 U261 (.IN1(new_block[16]), .IN2(n489), .IN3(new_block[48]), .IN4(n383), .IN5(
          n299), .Q(sboxw[16]));
   AO22X1 U262 (.IN1(new_block[112]), .IN2(n572), .IN3(new_block[80]), .IN4(n1315), .Q(
          n299));
   AO221X1 U263 (.IN1(new_block[15]), .IN2(n489), .IN3(new_block[47]), .IN4(n383), .IN5(
          n300), .Q(sboxw[15]));
   AO22X1 U264 (.IN1(new_block[111]), .IN2(n572), .IN3(new_block[79]), .IN4(n440), .Q(n300)
          );
   AO221X1 U265 (.IN1(new_block[14]), .IN2(n489), .IN3(new_block[46]), .IN4(n383), .IN5(
          n301), .Q(sboxw[14]));
   AO22X1 U266 (.IN1(new_block[110]), .IN2(n572), .IN3(new_block[78]), .IN4(n440), .Q(n301)
          );
   AO221X1 U267 (.IN1(new_block[13]), .IN2(n1316), .IN3(new_block[45]), .IN4(n383), .IN5(
          n302), .Q(sboxw[13]));
   AO22X1 U268 (.IN1(new_block[109]), .IN2(n572), .IN3(new_block[77]), .IN4(n1315), .Q(
          n302));
   AO221X1 U269 (.IN1(new_block[12]), .IN2(n489), .IN3(new_block[44]), .IN4(n383), .IN5(
          n303), .Q(sboxw[12]));
   AO22X1 U270 (.IN1(new_block[108]), .IN2(n572), .IN3(new_block[76]), .IN4(n440), .Q(n303)
          );
   AO221X1 U271 (.IN1(new_block[11]), .IN2(n489), .IN3(new_block[43]), .IN4(n383), .IN5(
          n304), .Q(sboxw[11]));
   AO22X1 U272 (.IN1(new_block[107]), .IN2(n572), .IN3(new_block[75]), .IN4(n440), .Q(n304)
          );
   AO221X1 U273 (.IN1(new_block[10]), .IN2(n489), .IN3(new_block[42]), .IN4(n383), .IN5(
          n305), .Q(sboxw[10]));
   AO22X1 U274 (.IN1(new_block[106]), .IN2(n572), .IN3(new_block[74]), .IN4(n440), .Q(n305)
          );
   AO221X1 U275 (.IN1(new_block[0]), .IN2(n1316), .IN3(new_block[32]), .IN4(n383), .IN5(
          n306), .Q(sboxw[0]));
   AO22X1 U276 (.IN1(new_block[96]), .IN2(n572), .IN3(new_block[64]), .IN4(n1315), .Q(n306)
          );
   AO221X1 U277 (.IN1(new_sboxw[31]), .IN2(n1265), .IN3(n592), .IN4(new_block[127]), .IN5(
          n312), .Q(n1117));
   AO22X1 U278 (.IN1(round_key[127]), .IN2(n313), .IN3(n314), .IN4(n1283), .Q(n312));
   AO222X1 U279 (.IN1(block[127]), .IN2(n966), .IN3(n1260), .IN4(n315), .IN5(n1254), .IN6(
          new_block[127]), .Q(n314));
   OAI222X1 U280 (.IN1(n315), .IN2(n316), .IN3(n1072), .IN4(new_block[127]), .IN5(n888), .
          IN6(block[127]), .QN(n313));
   XOR3X1 U281 (.IN1(new_block[47]), .IN2(n218), .IN3(n319), .Q(n315));
   XOR3X1 U282 (.IN1(new_block[87]), .IN2(new_block[86]), .IN3(n169), .Q(n319));
   AO221X1 U283 (.IN1(new_sboxw[30]), .IN2(n1265), .IN3(n579), .IN4(new_block[126]), .IN5(
          n320), .Q(n1118));
   AO22X1 U284 (.IN1(round_key[126]), .IN2(n321), .IN3(n322), .IN4(n1284), .Q(n320));
   AO222X1 U285 (.IN1(block[126]), .IN2(n897), .IN3(n433), .IN4(n323), .IN5(n1036), .IN6(
          new_block[126]), .Q(n322));
   OAI222X1 U286 (.IN1(n323), .IN2(n316), .IN3(n1084), .IN4(new_block[126]), .IN5(n876), .
          IN6(block[126]), .QN(n321));
   XNOR3X1 U287 (.IN1(new_block[46]), .IN2(new_block[125]), .IN3(n324), .Q(n323));
   XOR3X1 U288 (.IN1(new_block[86]), .IN2(new_block[85]), .IN3(n170), .Q(n324));
   AO221X1 U289 (.IN1(new_sboxw[29]), .IN2(n1265), .IN3(n579), .IN4(new_block[125]), .IN5(
          n325), .Q(n1119));
   AO22X1 U290 (.IN1(round_key[125]), .IN2(n326), .IN3(n327), .IN4(n1285), .Q(n325));
   AO222X1 U291 (.IN1(block[125]), .IN2(n840), .IN3(n1255), .IN4(n328), .IN5(n973), .IN6(
          new_block[125]), .Q(n327));
   OAI222X1 U292 (.IN1(n328), .IN2(n316), .IN3(n317), .IN4(new_block[125]), .IN5(n888), .
          IN6(block[125]), .QN(n326));
   XNOR3X1 U293 (.IN1(new_block[45]), .IN2(new_block[124]), .IN3(n329), .Q(n328));
   XOR3X1 U294 (.IN1(new_block[85]), .IN2(new_block[84]), .IN3(n171), .Q(n329));
   AO221X1 U295 (.IN1(new_sboxw[28]), .IN2(n1265), .IN3(n592), .IN4(new_block[124]), .IN5(
          n330), .Q(n1120));
   AO22X1 U296 (.IN1(round_key[124]), .IN2(n331), .IN3(n332), .IN4(n1286), .Q(n330));
   AO222X1 U297 (.IN1(block[124]), .IN2(n840), .IN3(n1255), .IN4(n333), .IN5(n403), .IN6(
          new_block[124]), .Q(n332));
   OAI222X1 U298 (.IN1(n333), .IN2(n316), .IN3(n317), .IN4(new_block[124]), .IN5(n888), .
          IN6(block[124]), .QN(n331));
   XNOR3X1 U299 (.IN1(n334), .IN2(n335), .IN3(n336), .Q(n333));
   XOR3X1 U300 (.IN1(new_block[84]), .IN2(n172), .IN3(new_block[44]), .Q(n336));
   AO221X1 U301 (.IN1(new_sboxw[27]), .IN2(n1265), .IN3(n579), .IN4(new_block[123]), .IN5(
          n337), .Q(n1121));
   AO22X1 U302 (.IN1(round_key[123]), .IN2(n338), .IN3(n339), .IN4(n1287), .Q(n337));
   AO222X1 U303 (.IN1(block[123]), .IN2(n777), .IN3(n433), .IN4(n340), .IN5(n973), .IN6(
          new_block[123]), .Q(n339));
   OAI222X1 U304 (.IN1(n340), .IN2(n316), .IN3(n317), .IN4(new_block[123]), .IN5(n876), .
          IN6(block[123]), .QN(n338));
   XNOR3X1 U305 (.IN1(n341), .IN2(n342), .IN3(n343), .Q(n340));
   XOR3X1 U306 (.IN1(new_block[83]), .IN2(new_block[43]), .IN3(n173), .Q(n343));
   AO221X1 U307 (.IN1(new_sboxw[26]), .IN2(n1265), .IN3(n592), .IN4(new_block[122]), .IN5(
          n344), .Q(n1122));
   AO22X1 U308 (.IN1(round_key[122]), .IN2(n345), .IN3(n346), .IN4(n1288), .Q(n344));
   AO222X1 U309 (.IN1(block[122]), .IN2(n390), .IN3(n1258), .IN4(n347), .IN5(n1066), .IN6(
          new_block[122]), .Q(n346));
   OAI222X1 U310 (.IN1(n347), .IN2(n1262), .IN3(n317), .IN4(new_block[122]), .IN5(n876), .
          IN6(block[122]), .QN(n345));
   XOR3X1 U311 (.IN1(new_block[2]), .IN2(n221), .IN3(n348), .Q(n347));
   XOR3X1 U312 (.IN1(new_block[82]), .IN2(new_block[81]), .IN3(n194), .Q(n348));
   AO221X1 U313 (.IN1(new_sboxw[25]), .IN2(n1265), .IN3(n579), .IN4(new_block[121]), .IN5(
          n349), .Q(n1123));
   AO22X1 U314 (.IN1(round_key[121]), .IN2(n350), .IN3(n351), .IN4(n1289), .Q(n349));
   AO222X1 U315 (.IN1(block[121]), .IN2(n966), .IN3(n1260), .IN4(n352), .IN5(n973), .IN6(
          new_block[121]), .Q(n351));
   OAI222X1 U316 (.IN1(n352), .IN2(n1263), .IN3(n317), .IN4(new_block[121]), .IN5(n888), .
          IN6(block[121]), .QN(n350));
   XNOR3X1 U317 (.IN1(n353), .IN2(n354), .IN3(n355), .Q(n352));
   XOR3X1 U318 (.IN1(new_block[81]), .IN2(n195), .IN3(new_block[1]), .Q(n355));
   AO221X1 U319 (.IN1(new_sboxw[24]), .IN2(n1265), .IN3(n592), .IN4(new_block[120]), .IN5(
          n356), .Q(n1124));
   AO22X1 U320 (.IN1(round_key[120]), .IN2(n357), .IN3(n358), .IN4(n1290), .Q(n356));
   AO222X1 U321 (.IN1(block[120]), .IN2(n897), .IN3(n1259), .IN4(n359), .IN5(n1113), .IN6(
          new_block[120]), .Q(n358));
   OAI222X1 U322 (.IN1(n359), .IN2(n1263), .IN3(n317), .IN4(new_block[120]), .IN5(n318), .
          IN6(block[120]), .QN(n357));
   XOR3X1 U323 (.IN1(n196), .IN2(new_block[127]), .IN3(n360), .Q(n359));
   XNOR2X1 U324 (.IN1(new_block[0]), .IN2(n353), .Q(n360));
   AO221X1 U325 (.IN1(n777), .IN2(n361), .IN3(n592), .IN4(new_block[119]), .IN5(n362), .Q(
          n1125));
   AO222X1 U326 (.IN1(new_sboxw[23]), .IN2(n1265), .IN3(n1254), .IN4(n363), .IN5(n1260), .
          IN6(n364), .Q(n362));
   XNOR3X1 U327 (.IN1(n365), .IN2(new_block[127]), .IN3(n366), .Q(n364));
   XOR3X1 U328 (.IN1(round_key[119]), .IN2(new_block[86]), .IN3(n169), .Q(n366));
   XOR2X1 U329 (.IN1(new_block[47]), .IN2(new_block[46]), .Q(n365));
   XOR2X1 U330 (.IN1(round_key[119]), .IN2(new_block[87]), .Q(n363));
   XOR2X1 U331 (.IN1(round_key[119]), .IN2(block[119]), .Q(n361));
   AO221X1 U332 (.IN1(n777), .IN2(n367), .IN3(n592), .IN4(new_block[118]), .IN5(n368), .Q(
          n1126));
   AO222X1 U333 (.IN1(new_sboxw[22]), .IN2(n1265), .IN3(n403), .IN4(n369), .IN5(n1258), .
          IN6(n370), .Q(n368));
   XOR3X1 U334 (.IN1(n371), .IN2(n218), .IN3(n372), .Q(n370));
   XOR3X1 U335 (.IN1(round_key[118]), .IN2(new_block[85]), .IN3(n170), .Q(n372));
   XOR2X1 U336 (.IN1(new_block[46]), .IN2(new_block[45]), .Q(n371));
   XOR2X1 U337 (.IN1(round_key[118]), .IN2(new_block[86]), .Q(n369));
   XOR2X1 U338 (.IN1(round_key[118]), .IN2(block[118]), .Q(n367));
   AO221X1 U339 (.IN1(n777), .IN2(n373), .IN3(n592), .IN4(new_block[117]), .IN5(n374), .Q(
          n1127));
   AO222X1 U340 (.IN1(new_sboxw[21]), .IN2(n1265), .IN3(n1036), .IN4(n375), .IN5(n433), .
          IN6(n376), .Q(n374));
   XOR3X1 U341 (.IN1(n377), .IN2(n219), .IN3(n378), .Q(n376));
   XOR3X1 U342 (.IN1(round_key[117]), .IN2(new_block[84]), .IN3(n171), .Q(n378));
   XOR2X1 U343 (.IN1(new_block[45]), .IN2(new_block[44]), .Q(n377));
   XOR2X1 U344 (.IN1(round_key[117]), .IN2(new_block[85]), .Q(n375));
   XOR2X1 U345 (.IN1(round_key[117]), .IN2(block[117]), .Q(n373));
   AO221X1 U346 (.IN1(n790), .IN2(n379), .IN3(n592), .IN4(new_block[116]), .IN5(n380), .Q(
          n1128));
   AO222X1 U347 (.IN1(new_sboxw[20]), .IN2(n1265), .IN3(n1254), .IN4(n381), .IN5(n1255), .
          IN6(n382), .Q(n380));
   XOR3X1 U349 (.IN1(n334), .IN2(new_block[124]), .IN3(n385), .Q(n384));
   XOR2X1 U350 (.IN1(new_block[83]), .IN2(new_block[87]), .Q(n334));
   XOR2X1 U352 (.IN1(round_key[116]), .IN2(new_block[84]), .Q(n381));
   XOR2X1 U353 (.IN1(round_key[116]), .IN2(block[116]), .Q(n379));
   AO221X1 U354 (.IN1(n777), .IN2(n386), .IN3(n592), .IN4(new_block[115]), .IN5(n387), .Q(
          n1129));
   AO222X1 U355 (.IN1(new_sboxw[19]), .IN2(n1265), .IN3(n1113), .IN4(n388), .IN5(n1260), .
          IN6(n389), .Q(n387));
   XOR3X1 U357 (.IN1(n341), .IN2(new_block[123]), .IN3(n392), .Q(n391));
   XOR2X1 U358 (.IN1(new_block[82]), .IN2(new_block[87]), .Q(n341));
   XOR2X1 U360 (.IN1(round_key[115]), .IN2(new_block[83]), .Q(n388));
   XOR2X1 U361 (.IN1(round_key[115]), .IN2(block[115]), .Q(n386));
   AO221X1 U362 (.IN1(n790), .IN2(n393), .IN3(n592), .IN4(new_block[114]), .IN5(n394), .Q(
          n1130));
   AO222X1 U363 (.IN1(new_sboxw[18]), .IN2(n1266), .IN3(n973), .IN4(n395), .IN5(n1261), .
          IN6(n396), .Q(n394));
   XOR3X1 U364 (.IN1(n397), .IN2(n220), .IN3(n398), .Q(n396));
   XOR3X1 U365 (.IN1(round_key[114]), .IN2(new_block[81]), .IN3(n194), .Q(n398));
   XOR2X1 U366 (.IN1(new_block[41]), .IN2(new_block[2]), .Q(n397));
   XOR2X1 U367 (.IN1(round_key[114]), .IN2(new_block[82]), .Q(n395));
   XOR2X1 U368 (.IN1(round_key[114]), .IN2(block[114]), .Q(n393));
   AO221X1 U369 (.IN1(n820), .IN2(n399), .IN3(n592), .IN4(new_block[113]), .IN5(n400), .Q(
          n1131));
   AO222X1 U370 (.IN1(new_sboxw[17]), .IN2(n1266), .IN3(n1023), .IN4(n401), .IN5(n1260), .
          IN6(n402), .Q(n400));
   XOR3X1 U372 (.IN1(n353), .IN2(new_block[121]), .IN3(n405), .Q(n404));
   XOR2X1 U373 (.IN1(new_block[80]), .IN2(new_block[87]), .Q(n353));
   XOR2X1 U375 (.IN1(round_key[113]), .IN2(new_block[81]), .Q(n401));
   XOR2X1 U376 (.IN1(round_key[113]), .IN2(block[113]), .Q(n399));
   AO221X1 U377 (.IN1(n827), .IN2(n406), .IN3(n592), .IN4(new_block[112]), .IN5(n407), .Q(
          n1132));
   AO222X1 U378 (.IN1(new_sboxw[16]), .IN2(n1266), .IN3(n1066), .IN4(n408), .IN5(n1257), .
          IN6(n409), .Q(n407));
   XNOR3X1 U379 (.IN1(n405), .IN2(new_block[0]), .IN3(n410), .Q(n409));
   XOR2X1 U381 (.IN1(round_key[112]), .IN2(new_block[80]), .Q(n408));
   XOR2X1 U382 (.IN1(round_key[112]), .IN2(block[112]), .Q(n406));
   AO221X1 U383 (.IN1(n870), .IN2(n411), .IN3(n592), .IN4(new_block[111]), .IN5(n412), .Q(
          n1133));
   AO222X1 U384 (.IN1(new_sboxw[15]), .IN2(n1266), .IN3(n1113), .IN4(n413), .IN5(n433), .
          IN6(n414), .Q(n412));
   XNOR3X1 U385 (.IN1(n415), .IN2(new_block[127]), .IN3(n416), .Q(n414));
   XOR3X1 U386 (.IN1(round_key[111]), .IN2(new_block[87]), .IN3(n169), .Q(n416));
   XOR2X1 U387 (.IN1(new_block[6]), .IN2(new_block[46]), .Q(n415));
   XOR2X1 U388 (.IN1(round_key[111]), .IN2(new_block[47]), .Q(n413));
   XOR2X1 U389 (.IN1(round_key[111]), .IN2(block[111]), .Q(n411));
   AO221X1 U390 (.IN1(n870), .IN2(n417), .IN3(n592), .IN4(new_block[110]), .IN5(n418), .Q(
          n1134));
   AO222X1 U391 (.IN1(new_sboxw[14]), .IN2(n1266), .IN3(n1036), .IN4(n419), .IN5(n1258), .
          IN6(n420), .Q(n418));
   XOR3X1 U392 (.IN1(n421), .IN2(n218), .IN3(n422), .Q(n420));
   XOR3X1 U393 (.IN1(round_key[110]), .IN2(new_block[86]), .IN3(n170), .Q(n422));
   XOR2X1 U394 (.IN1(new_block[5]), .IN2(new_block[45]), .Q(n421));
   XOR2X1 U395 (.IN1(round_key[110]), .IN2(new_block[46]), .Q(n419));
   XOR2X1 U396 (.IN1(round_key[110]), .IN2(block[110]), .Q(n417));
   AO221X1 U397 (.IN1(n790), .IN2(n423), .IN3(n592), .IN4(new_block[109]), .IN5(n424), .Q(
          n1135));
   AO222X1 U398 (.IN1(new_sboxw[13]), .IN2(n1266), .IN3(n986), .IN4(n425), .IN5(n1264), .
          IN6(n426), .Q(n424));
   XOR3X1 U399 (.IN1(n427), .IN2(n219), .IN3(n428), .Q(n426));
   XOR3X1 U400 (.IN1(round_key[109]), .IN2(new_block[85]), .IN3(n171), .Q(n428));
   XOR2X1 U401 (.IN1(new_block[4]), .IN2(new_block[44]), .Q(n427));
   XOR2X1 U402 (.IN1(round_key[109]), .IN2(new_block[45]), .Q(n425));
   XOR2X1 U403 (.IN1(round_key[109]), .IN2(block[109]), .Q(n423));
   AO221X1 U404 (.IN1(n840), .IN2(n429), .IN3(n592), .IN4(new_block[108]), .IN5(n430), .Q(
          n1136));
   AO222X1 U405 (.IN1(new_sboxw[12]), .IN2(n1266), .IN3(n973), .IN4(n431), .IN5(n1259), .
          IN6(n432), .Q(n430));
   XNOR3X1 U407 (.IN1(n385), .IN2(new_block[124]), .IN3(n435), .Q(n434));
   XOR2X1 U408 (.IN1(n193), .IN2(n192), .Q(n385));
   XOR2X1 U410 (.IN1(round_key[108]), .IN2(new_block[44]), .Q(n431));
   XOR2X1 U411 (.IN1(round_key[108]), .IN2(block[108]), .Q(n429));
   AO221X1 U412 (.IN1(n820), .IN2(n436), .IN3(n579), .IN4(new_block[107]), .IN5(n437), .Q(
          n1137));
   AO222X1 U413 (.IN1(new_sboxw[11]), .IN2(n1266), .IN3(n1036), .IN4(n438), .IN5(n433), .
          IN6(n439), .Q(n437));
   XNOR3X1 U415 (.IN1(n392), .IN2(new_block[123]), .IN3(n442), .Q(n441));
   XOR2X1 U416 (.IN1(n194), .IN2(n192), .Q(n392));
   XOR2X1 U418 (.IN1(round_key[107]), .IN2(new_block[43]), .Q(n438));
   XOR2X1 U419 (.IN1(round_key[107]), .IN2(block[107]), .Q(n436));
   AO221X1 U420 (.IN1(n827), .IN2(n443), .IN3(n579), .IN4(new_block[106]), .IN5(n444), .Q(
          n1138));
   AO222X1 U421 (.IN1(new_sboxw[10]), .IN2(n1266), .IN3(n1066), .IN4(n445), .IN5(n1264), .
          IN6(n446), .Q(n444));
   XOR3X1 U422 (.IN1(n447), .IN2(n220), .IN3(n448), .Q(n446));
   XOR3X1 U423 (.IN1(round_key[106]), .IN2(new_block[82]), .IN3(n195), .Q(n448));
   XOR2X1 U424 (.IN1(new_block[2]), .IN2(new_block[1]), .Q(n447));
   XOR2X1 U425 (.IN1(round_key[106]), .IN2(new_block[42]), .Q(n445));
   XOR2X1 U426 (.IN1(round_key[106]), .IN2(block[106]), .Q(n443));
   AO221X1 U427 (.IN1(n897), .IN2(n449), .IN3(n579), .IN4(new_block[105]), .IN5(n450), .Q(
          n1139));
   AO222X1 U428 (.IN1(new_sboxw[9]), .IN2(n1266), .IN3(n1016), .IN4(n451), .IN5(n1257), .
          IN6(n452), .Q(n450));
   XOR3X1 U430 (.IN1(n405), .IN2(n221), .IN3(n455), .Q(n454));
   XOR2X1 U431 (.IN1(n196), .IN2(n192), .Q(n405));
   XOR2X1 U433 (.IN1(round_key[105]), .IN2(new_block[41]), .Q(n451));
   XOR2X1 U434 (.IN1(round_key[105]), .IN2(block[105]), .Q(n449));
   AO221X1 U435 (.IN1(n820), .IN2(n456), .IN3(n579), .IN4(new_block[104]), .IN5(n457), .Q(
          n1140));
   AO222X1 U436 (.IN1(new_sboxw[8]), .IN2(n1266), .IN3(n1023), .IN4(n458), .IN5(n1261), .
          IN6(n459), .Q(n457));
   XOR3X1 U437 (.IN1(n455), .IN2(new_block[120]), .IN3(n460), .Q(n459));
   XOR3X1 U438 (.IN1(round_key[104]), .IN2(new_block[80]), .IN3(n192), .Q(n460));
   XOR2X1 U439 (.IN1(round_key[104]), .IN2(new_block[40]), .Q(n458));
   XOR2X1 U440 (.IN1(round_key[104]), .IN2(block[104]), .Q(n456));
   AO221X1 U441 (.IN1(n820), .IN2(n461), .IN3(n579), .IN4(new_block[103]), .IN5(n462), .Q(
          n1141));
   AO222X1 U442 (.IN1(new_sboxw[7]), .IN2(n1266), .IN3(n1066), .IN4(n463), .IN5(n1256), .
          IN6(n464), .Q(n462));
   XOR3X1 U443 (.IN1(n465), .IN2(n218), .IN3(n466), .Q(n464));
   XOR3X1 U444 (.IN1(round_key[103]), .IN2(new_block[87]), .IN3(n170), .Q(n466));
   XOR2X1 U445 (.IN1(new_block[47]), .IN2(new_block[127]), .Q(n465));
   XOR2X1 U446 (.IN1(round_key[103]), .IN2(new_block[7]), .Q(n463));
   XOR2X1 U447 (.IN1(round_key[103]), .IN2(block[103]), .Q(n461));
   AO221X1 U448 (.IN1(n827), .IN2(n467), .IN3(n579), .IN4(new_block[102]), .IN5(n468), .Q(
          n1142));
   AO222X1 U449 (.IN1(new_sboxw[6]), .IN2(n1266), .IN3(n1016), .IN4(n469), .IN5(n1259), .
          IN6(n470), .Q(n468));
   XOR3X1 U450 (.IN1(n471), .IN2(n219), .IN3(n472), .Q(n470));
   XOR3X1 U451 (.IN1(round_key[102]), .IN2(new_block[86]), .IN3(n171), .Q(n472));
   XOR2X1 U452 (.IN1(new_block[46]), .IN2(new_block[126]), .Q(n471));
   XOR2X1 U453 (.IN1(round_key[102]), .IN2(new_block[6]), .Q(n469));
   XOR2X1 U454 (.IN1(round_key[102]), .IN2(block[102]), .Q(n467));
   AO221X1 U455 (.IN1(n870), .IN2(n473), .IN3(n579), .IN4(new_block[101]), .IN5(n474), .Q(
          n1143));
   AO222X1 U456 (.IN1(new_sboxw[5]), .IN2(n1266), .IN3(n986), .IN4(n475), .IN5(n433), .IN6(
          n476), .Q(n474));
   XNOR3X1 U457 (.IN1(n477), .IN2(new_block[124]), .IN3(n478), .Q(n476));
   XOR3X1 U458 (.IN1(round_key[101]), .IN2(new_block[85]), .IN3(n172), .Q(n478));
   XOR2X1 U459 (.IN1(new_block[45]), .IN2(new_block[125]), .Q(n477));
   XOR2X1 U460 (.IN1(round_key[101]), .IN2(new_block[5]), .Q(n475));
   XOR2X1 U461 (.IN1(round_key[101]), .IN2(block[101]), .Q(n473));
   AO221X1 U462 (.IN1(n790), .IN2(n479), .IN3(n579), .IN4(new_block[100]), .IN5(n480), .Q(
          n1144));
   AO222X1 U463 (.IN1(new_sboxw[4]), .IN2(n1265), .IN3(n1023), .IN4(n481), .IN5(n1260), .
          IN6(n482), .Q(n480));
   XNOR3X1 U465 (.IN1(n335), .IN2(new_block[124]), .IN3(n435), .Q(n484));
   XOR2X1 U466 (.IN1(n173), .IN2(new_block[7]), .Q(n435));
   XOR2X1 U467 (.IN1(new_block[123]), .IN2(new_block[127]), .Q(n335));
   XOR2X1 U469 (.IN1(round_key[100]), .IN2(new_block[4]), .Q(n481));
   XOR2X1 U470 (.IN1(round_key[100]), .IN2(block[100]), .Q(n479));
   AO221X1 U471 (.IN1(n840), .IN2(n485), .IN3(n579), .IN4(new_block[99]), .IN5(n486), .Q(
          n1145));
   AO222X1 U472 (.IN1(new_sboxw[3]), .IN2(n1265), .IN3(n986), .IN4(n487), .IN5(n1261), .
          IN6(n488), .Q(n486));
   XNOR3X1 U474 (.IN1(n342), .IN2(new_block[123]), .IN3(n442), .Q(n490));
   XOR2X1 U475 (.IN1(n174), .IN2(new_block[7]), .Q(n442));
   XOR2X1 U476 (.IN1(new_block[122]), .IN2(new_block[127]), .Q(n342));
   XOR2X1 U478 (.IN1(round_key[99]), .IN2(new_block[3]), .Q(n487));
   XOR2X1 U479 (.IN1(round_key[99]), .IN2(block[99]), .Q(n485));
   AO221X1 U480 (.IN1(n790), .IN2(n491), .IN3(n579), .IN4(new_block[98]), .IN5(n492), .Q(
          n1146));
   AO222X1 U481 (.IN1(new_sboxw[2]), .IN2(n1266), .IN3(n1254), .IN4(n493), .IN5(n1257), .
          IN6(n494), .Q(n492));
   XOR3X1 U482 (.IN1(n495), .IN2(n221), .IN3(n496), .Q(n494));
   XOR3X1 U483 (.IN1(round_key[98]), .IN2(new_block[82]), .IN3(n194), .Q(n496));
   XOR2X1 U484 (.IN1(new_block[1]), .IN2(new_block[122]), .Q(n495));
   XOR2X1 U485 (.IN1(round_key[98]), .IN2(new_block[2]), .Q(n493));
   XOR2X1 U486 (.IN1(round_key[98]), .IN2(block[98]), .Q(n491));
   AO221X1 U487 (.IN1(n897), .IN2(n497), .IN3(n579), .IN4(new_block[97]), .IN5(n498), .Q(
          n1147));
   AO222X1 U488 (.IN1(new_sboxw[1]), .IN2(n1265), .IN3(n1113), .IN4(n499), .IN5(n1261), .
          IN6(n500), .Q(n498));
   XOR3X1 U490 (.IN1(n354), .IN2(n221), .IN3(n455), .Q(n502));
   XOR2X1 U491 (.IN1(new_block[0]), .IN2(n169), .Q(n455));
   XOR2X1 U493 (.IN1(round_key[97]), .IN2(new_block[1]), .Q(n499));
   XOR2X1 U494 (.IN1(round_key[97]), .IN2(block[97]), .Q(n497));
   AO221X1 U495 (.IN1(n701), .IN2(new_sboxw[31]), .IN3(n483), .IN4(new_block[95]), .IN5(
          n504), .Q(n1148));
   AO22X1 U496 (.IN1(round_key[95]), .IN2(n505), .IN3(n506), .IN4(n1291), .Q(n504));
   AO222X1 U497 (.IN1(block[95]), .IN2(n777), .IN3(n1256), .IN4(n507), .IN5(n986), .IN6(
          new_block[95]), .Q(n506));
   OAI222X1 U498 (.IN1(n507), .IN2(n316), .IN3(n317), .IN4(new_block[95]), .IN5(n888), .
          IN6(block[95]), .QN(n505));
   XOR3X1 U499 (.IN1(new_block[15]), .IN2(n236), .IN3(n508), .Q(n507));
   XOR3X1 U500 (.IN1(new_block[94]), .IN2(new_block[55]), .IN3(n186), .Q(n508));
   AO221X1 U501 (.IN1(n701), .IN2(new_sboxw[30]), .IN3(n453), .IN4(new_block[94]), .IN5(
          n509), .Q(n1149));
   AO22X1 U502 (.IN1(round_key[94]), .IN2(n510), .IN3(n511), .IN4(n1292), .Q(n509));
   AO222X1 U503 (.IN1(block[94]), .IN2(n897), .IN3(n1257), .IN4(n512), .IN5(n1113), .IN6(
          new_block[94]), .Q(n511));
   OAI222X1 U504 (.IN1(n512), .IN2(n1262), .IN3(n1072), .IN4(new_block[94]), .IN5(n876), .
          IN6(block[94]), .QN(n510));
   XNOR3X1 U505 (.IN1(new_block[14]), .IN2(new_block[102]), .IN3(n513), .Q(n512));
   XOR3X1 U506 (.IN1(new_block[93]), .IN2(new_block[54]), .IN3(n187), .Q(n513));
   AO221X1 U507 (.IN1(n701), .IN2(new_sboxw[29]), .IN3(n483), .IN4(new_block[93]), .IN5(
          n514), .Q(n1150));
   AO22X1 U508 (.IN1(round_key[93]), .IN2(n515), .IN3(n516), .IN4(n1293), .Q(n514));
   AO222X1 U509 (.IN1(block[93]), .IN2(n870), .IN3(n1257), .IN4(n517), .IN5(n1023), .IN6(
          new_block[93]), .Q(n516));
   OAI222X1 U510 (.IN1(n517), .IN2(n1262), .IN3(n1084), .IN4(new_block[93]), .IN5(n888), .
          IN6(block[93]), .QN(n515));
   XNOR3X1 U511 (.IN1(new_block[13]), .IN2(new_block[101]), .IN3(n518), .Q(n517));
   XOR3X1 U512 (.IN1(new_block[92]), .IN2(new_block[53]), .IN3(n188), .Q(n518));
   AO221X1 U513 (.IN1(n701), .IN2(new_sboxw[28]), .IN3(n453), .IN4(new_block[92]), .IN5(
          n519), .Q(n1151));
   AO22X1 U514 (.IN1(round_key[92]), .IN2(n520), .IN3(n521), .IN4(n1294), .Q(n519));
   AO222X1 U515 (.IN1(block[92]), .IN2(n820), .IN3(n1264), .IN4(n522), .IN5(n1066), .IN6(
          new_block[92]), .Q(n521));
   OAI222X1 U516 (.IN1(n522), .IN2(n1263), .IN3(n1072), .IN4(new_block[92]), .IN5(n318), .
          IN6(block[92]), .QN(n520));
   XNOR3X1 U517 (.IN1(n523), .IN2(n524), .IN3(n525), .Q(n522));
   XOR3X1 U518 (.IN1(new_block[52]), .IN2(new_block[12]), .IN3(n239), .Q(n525));
   AO221X1 U519 (.IN1(n701), .IN2(new_sboxw[27]), .IN3(n483), .IN4(new_block[91]), .IN5(
          n526), .Q(n1152));
   AO22X1 U520 (.IN1(round_key[91]), .IN2(n527), .IN3(n528), .IN4(n1295), .Q(n526));
   AO222X1 U521 (.IN1(block[91]), .IN2(n790), .IN3(n1258), .IN4(n529), .IN5(n1254), .IN6(
          new_block[91]), .Q(n528));
   OAI222X1 U522 (.IN1(n529), .IN2(n316), .IN3(n317), .IN4(new_block[91]), .IN5(n888), .
          IN6(block[91]), .QN(n527));
   XNOR3X1 U523 (.IN1(n530), .IN2(n531), .IN3(n532), .Q(n529));
   XOR3X1 U524 (.IN1(new_block[99]), .IN2(new_block[51]), .IN3(n167), .Q(n532));
   AO221X1 U525 (.IN1(n701), .IN2(new_sboxw[26]), .IN3(n453), .IN4(new_block[90]), .IN5(
          n533), .Q(n1153));
   AO22X1 U526 (.IN1(round_key[90]), .IN2(n534), .IN3(n535), .IN4(n1296), .Q(n533));
   AO222X1 U527 (.IN1(block[90]), .IN2(n390), .IN3(n1264), .IN4(n536), .IN5(n1023), .IN6(
          new_block[90]), .Q(n535));
   OAI222X1 U528 (.IN1(n536), .IN2(n1262), .IN3(n1072), .IN4(new_block[90]), .IN5(n876), .
          IN6(block[90]), .QN(n534));
   XOR3X1 U529 (.IN1(new_block[49]), .IN2(n168), .IN3(n537), .Q(n536));
   XOR3X1 U530 (.IN1(new_block[98]), .IN2(new_block[89]), .IN3(n190), .Q(n537));
   AO221X1 U531 (.IN1(n701), .IN2(new_sboxw[25]), .IN3(n483), .IN4(new_block[89]), .IN5(
          n538), .Q(n1154));
   AO22X1 U532 (.IN1(round_key[89]), .IN2(n539), .IN3(n540), .IN4(n1297), .Q(n538));
   AO222X1 U533 (.IN1(block[89]), .IN2(n790), .IN3(n433), .IN4(n541), .IN5(n1113), .IN6(
          new_block[89]), .Q(n540));
   OAI222X1 U534 (.IN1(n541), .IN2(n1263), .IN3(n1084), .IN4(new_block[89]), .IN5(n876), .
          IN6(block[89]), .QN(n539));
   XNOR3X1 U535 (.IN1(n542), .IN2(n543), .IN3(n544), .Q(n541));
   XOR3X1 U536 (.IN1(new_block[9]), .IN2(new_block[97]), .IN3(n191), .Q(n544));
   AO221X1 U537 (.IN1(n701), .IN2(new_sboxw[24]), .IN3(n453), .IN4(new_block[88]), .IN5(
          n545), .Q(n1155));
   AO22X1 U538 (.IN1(round_key[88]), .IN2(n546), .IN3(n547), .IN4(n1298), .Q(n545));
   AO222X1 U539 (.IN1(block[88]), .IN2(n840), .IN3(n433), .IN4(n548), .IN5(n403), .IN6(
          new_block[88]), .Q(n547));
   OAI222X1 U540 (.IN1(n548), .IN2(n1263), .IN3(n1072), .IN4(new_block[88]), .IN5(n876), .
          IN6(block[88]), .QN(n546));
   XNOR3X1 U541 (.IN1(new_block[96]), .IN2(new_block[95]), .IN3(n549), .Q(n548));
   XNOR2X1 U542 (.IN1(new_block[8]), .IN2(n542), .Q(n549));
   AO221X1 U543 (.IN1(n390), .IN2(n550), .IN3(n483), .IN4(new_block[87]), .IN5(n551), .Q(
          n1156));
   AO222X1 U544 (.IN1(n701), .IN2(new_sboxw[23]), .IN3(n1066), .IN4(n552), .IN5(n1255), .
          IN6(n553), .Q(n551));
   XOR3X1 U545 (.IN1(n554), .IN2(n236), .IN3(n555), .Q(n553));
   XOR3X1 U546 (.IN1(round_key[87]), .IN2(new_block[95]), .IN3(n186), .Q(n555));
   XOR2X1 U547 (.IN1(new_block[15]), .IN2(new_block[14]), .Q(n554));
   XOR2X1 U548 (.IN1(round_key[87]), .IN2(new_block[55]), .Q(n552));
   XOR2X1 U549 (.IN1(round_key[87]), .IN2(block[87]), .Q(n550));
   AO221X1 U550 (.IN1(n840), .IN2(n556), .IN3(n483), .IN4(new_block[86]), .IN5(n557), .Q(
          n1157));
   AO222X1 U551 (.IN1(n701), .IN2(new_sboxw[22]), .IN3(n1023), .IN4(n558), .IN5(n1255), .
          IN6(n559), .Q(n557));
   XOR3X1 U552 (.IN1(n560), .IN2(n237), .IN3(n561), .Q(n559));
   XOR3X1 U553 (.IN1(round_key[86]), .IN2(new_block[94]), .IN3(n187), .Q(n561));
   XOR2X1 U554 (.IN1(new_block[14]), .IN2(new_block[13]), .Q(n560));
   XOR2X1 U555 (.IN1(round_key[86]), .IN2(new_block[54]), .Q(n558));
   XOR2X1 U556 (.IN1(round_key[86]), .IN2(block[86]), .Q(n556));
   AO221X1 U557 (.IN1(n966), .IN2(n562), .IN3(n483), .IN4(new_block[85]), .IN5(n563), .Q(
          n1158));
   AO222X1 U558 (.IN1(n701), .IN2(new_sboxw[21]), .IN3(n403), .IN4(n564), .IN5(n1261), .
          IN6(n565), .Q(n563));
   XOR3X1 U559 (.IN1(n566), .IN2(n238), .IN3(n567), .Q(n565));
   XOR3X1 U560 (.IN1(round_key[85]), .IN2(new_block[93]), .IN3(n188), .Q(n567));
   XOR2X1 U561 (.IN1(new_block[13]), .IN2(new_block[12]), .Q(n566));
   XOR2X1 U562 (.IN1(round_key[85]), .IN2(new_block[53]), .Q(n564));
   XOR2X1 U563 (.IN1(round_key[85]), .IN2(block[85]), .Q(n562));
   AO221X1 U564 (.IN1(n390), .IN2(n568), .IN3(n483), .IN4(new_block[84]), .IN5(n569), .Q(
          n1159));
   AO222X1 U565 (.IN1(n701), .IN2(new_sboxw[20]), .IN3(n1036), .IN4(n570), .IN5(n1260), .
          IN6(n571), .Q(n569));
   XOR3X1 U567 (.IN1(n523), .IN2(new_block[100]), .IN3(n574), .Q(n573));
   XOR2X1 U568 (.IN1(new_block[51]), .IN2(new_block[55]), .Q(n523));
   XOR2X1 U570 (.IN1(round_key[84]), .IN2(new_block[52]), .Q(n570));
   XOR2X1 U571 (.IN1(round_key[84]), .IN2(block[84]), .Q(n568));
   AO221X1 U572 (.IN1(n870), .IN2(n575), .IN3(n483), .IN4(new_block[83]), .IN5(n576), .Q(
          n1160));
   AO222X1 U573 (.IN1(n701), .IN2(new_sboxw[19]), .IN3(n1036), .IN4(n577), .IN5(n1261), .
          IN6(n578), .Q(n576));
   XOR3X1 U575 (.IN1(n530), .IN2(new_block[11]), .IN3(n581), .Q(n580));
   XOR2X1 U576 (.IN1(new_block[50]), .IN2(new_block[55]), .Q(n530));
   XOR2X1 U578 (.IN1(round_key[83]), .IN2(new_block[51]), .Q(n577));
   XOR2X1 U579 (.IN1(round_key[83]), .IN2(block[83]), .Q(n575));
   AO221X1 U580 (.IN1(n840), .IN2(n582), .IN3(n483), .IN4(new_block[82]), .IN5(n583), .Q(
          n1161));
   AO222X1 U581 (.IN1(n770), .IN2(new_sboxw[18]), .IN3(n1113), .IN4(n584), .IN5(n1256), .
          IN6(n585), .Q(n583));
   XOR3X1 U582 (.IN1(n586), .IN2(n168), .IN3(n587), .Q(n585));
   XOR3X1 U583 (.IN1(round_key[82]), .IN2(new_block[9]), .IN3(n241), .Q(n587));
   XOR2X1 U584 (.IN1(new_block[90]), .IN2(new_block[49]), .Q(n586));
   XOR2X1 U585 (.IN1(round_key[82]), .IN2(new_block[50]), .Q(n584));
   XOR2X1 U586 (.IN1(round_key[82]), .IN2(block[82]), .Q(n582));
   AO221X1 U587 (.IN1(n777), .IN2(n588), .IN3(n483), .IN4(new_block[81]), .IN5(n589), .Q(
          n1162));
   AO222X1 U588 (.IN1(n770), .IN2(new_sboxw[17]), .IN3(n1036), .IN4(n590), .IN5(n1256), .
          IN6(n591), .Q(n589));
   XOR3X1 U590 (.IN1(n542), .IN2(new_block[89]), .IN3(n594), .Q(n593));
   XOR2X1 U591 (.IN1(new_block[48]), .IN2(new_block[55]), .Q(n542));
   XOR2X1 U593 (.IN1(round_key[81]), .IN2(new_block[49]), .Q(n590));
   XOR2X1 U594 (.IN1(round_key[81]), .IN2(block[81]), .Q(n588));
   AO221X1 U595 (.IN1(n790), .IN2(n595), .IN3(n483), .IN4(new_block[80]), .IN5(n596), .Q(
          n1163));
   AO222X1 U596 (.IN1(n770), .IN2(new_sboxw[16]), .IN3(n1113), .IN4(n597), .IN5(n1259), .
          IN6(n598), .Q(n596));
   XOR3X1 U597 (.IN1(n594), .IN2(n185), .IN3(n599), .Q(n598));
   XNOR3X1 U598 (.IN1(round_key[80]), .IN2(new_block[96]), .IN3(new_block[88]), .Q(n599)
          );
   XOR2X1 U599 (.IN1(round_key[80]), .IN2(new_block[48]), .Q(n597));
   XOR2X1 U600 (.IN1(round_key[80]), .IN2(block[80]), .Q(n595));
   AO221X1 U601 (.IN1(n777), .IN2(n600), .IN3(n483), .IN4(new_block[79]), .IN5(n601), .Q(
          n1164));
   AO222X1 U602 (.IN1(n770), .IN2(new_sboxw[15]), .IN3(n1016), .IN4(n602), .IN5(n1261), .
          IN6(n603), .Q(n601));
   XOR3X1 U603 (.IN1(n604), .IN2(n237), .IN3(n605), .Q(n603));
   XOR3X1 U604 (.IN1(round_key[79]), .IN2(new_block[95]), .IN3(n185), .Q(n605));
   XOR2X1 U605 (.IN1(new_block[14]), .IN2(new_block[103]), .Q(n604));
   XOR2X1 U606 (.IN1(round_key[79]), .IN2(new_block[15]), .Q(n602));
   XOR2X1 U607 (.IN1(round_key[79]), .IN2(block[79]), .Q(n600));
   AO221X1 U608 (.IN1(n390), .IN2(n606), .IN3(n483), .IN4(new_block[78]), .IN5(n607), .Q(
          n1165));
   AO222X1 U609 (.IN1(n770), .IN2(new_sboxw[14]), .IN3(n1066), .IN4(n608), .IN5(n1258), .
          IN6(n609), .Q(n607));
   XOR3X1 U610 (.IN1(n610), .IN2(n238), .IN3(n611), .Q(n609));
   XOR3X1 U611 (.IN1(round_key[78]), .IN2(new_block[94]), .IN3(n186), .Q(n611));
   XOR2X1 U612 (.IN1(new_block[13]), .IN2(new_block[102]), .Q(n610));
   XOR2X1 U613 (.IN1(round_key[78]), .IN2(new_block[14]), .Q(n608));
   XOR2X1 U614 (.IN1(round_key[78]), .IN2(block[78]), .Q(n606));
   AO221X1 U615 (.IN1(n827), .IN2(n612), .IN3(n483), .IN4(new_block[77]), .IN5(n613), .Q(
          n1166));
   AO222X1 U616 (.IN1(n770), .IN2(new_sboxw[13]), .IN3(n1066), .IN4(n614), .IN5(n1256), .
          IN6(n615), .Q(n613));
   XOR3X1 U617 (.IN1(n616), .IN2(n239), .IN3(n617), .Q(n615));
   XOR3X1 U618 (.IN1(round_key[77]), .IN2(new_block[93]), .IN3(n187), .Q(n617));
   XOR2X1 U619 (.IN1(new_block[12]), .IN2(new_block[101]), .Q(n616));
   XOR2X1 U620 (.IN1(round_key[77]), .IN2(new_block[13]), .Q(n614));
   XOR2X1 U621 (.IN1(round_key[77]), .IN2(block[77]), .Q(n612));
   AO221X1 U622 (.IN1(n777), .IN2(n618), .IN3(n483), .IN4(new_block[76]), .IN5(n619), .Q(
          n1167));
   AO222X1 U623 (.IN1(n770), .IN2(new_sboxw[12]), .IN3(n1016), .IN4(n620), .IN5(n1257), .
          IN6(n621), .Q(n619));
   XOR3X1 U625 (.IN1(n574), .IN2(n239), .IN3(n624), .Q(n623));
   XOR2X1 U626 (.IN1(n167), .IN2(n166), .Q(n574));
   XOR2X1 U628 (.IN1(round_key[76]), .IN2(new_block[12]), .Q(n620));
   XOR2X1 U629 (.IN1(round_key[76]), .IN2(block[76]), .Q(n618));
   AO221X1 U630 (.IN1(n790), .IN2(n625), .IN3(n453), .IN4(new_block[75]), .IN5(n626), .Q(
          n1168));
   AO222X1 U631 (.IN1(n770), .IN2(new_sboxw[11]), .IN3(n1023), .IN4(n627), .IN5(n433), .
          IN6(n628), .Q(n626));
   XOR3X1 U633 (.IN1(n581), .IN2(n189), .IN3(n631), .Q(n630));
   XOR2X1 U634 (.IN1(n168), .IN2(n166), .Q(n581));
   XOR2X1 U636 (.IN1(round_key[75]), .IN2(new_block[11]), .Q(n627));
   XOR2X1 U637 (.IN1(round_key[75]), .IN2(block[75]), .Q(n625));
   AO221X1 U638 (.IN1(n820), .IN2(n632), .IN3(n453), .IN4(new_block[74]), .IN5(n633), .Q(
          n1169));
   AO222X1 U639 (.IN1(n770), .IN2(new_sboxw[10]), .IN3(n1254), .IN4(n634), .IN5(n1255), .
          IN6(n635), .Q(n633));
   XOR3X1 U640 (.IN1(n636), .IN2(n190), .IN3(n637), .Q(n635));
   XOR3X1 U641 (.IN1(round_key[74]), .IN2(new_block[9]), .IN3(n241), .Q(n637));
   XOR2X1 U642 (.IN1(new_block[97]), .IN2(new_block[90]), .Q(n636));
   XOR2X1 U643 (.IN1(round_key[74]), .IN2(new_block[10]), .Q(n634));
   XOR2X1 U644 (.IN1(round_key[74]), .IN2(block[74]), .Q(n632));
   AO221X1 U645 (.IN1(n870), .IN2(n638), .IN3(n453), .IN4(new_block[73]), .IN5(n639), .Q(
          n1170));
   AO222X1 U646 (.IN1(n770), .IN2(new_sboxw[9]), .IN3(n1113), .IN4(n640), .IN5(n1256), .
          IN6(n641), .Q(n639));
   XOR3X1 U648 (.IN1(n594), .IN2(n191), .IN3(n644), .Q(n643));
   XOR2X1 U649 (.IN1(new_block[8]), .IN2(new_block[15]), .Q(n594));
   XOR2X1 U651 (.IN1(round_key[73]), .IN2(new_block[9]), .Q(n640));
   XOR2X1 U652 (.IN1(round_key[73]), .IN2(block[73]), .Q(n638));
   AO221X1 U653 (.IN1(n827), .IN2(n645), .IN3(n453), .IN4(new_block[72]), .IN5(n646), .Q(
          n1171));
   AO222X1 U654 (.IN1(n770), .IN2(new_sboxw[8]), .IN3(n1066), .IN4(n647), .IN5(n1260), .
          IN6(n648), .Q(n646));
   XOR3X1 U655 (.IN1(n644), .IN2(new_block[15]), .IN3(n649), .Q(n648));
   XNOR3X1 U656 (.IN1(round_key[72]), .IN2(new_block[88]), .IN3(new_block[48]), .Q(n649)
          );
   XOR2X1 U657 (.IN1(round_key[72]), .IN2(new_block[8]), .Q(n647));
   XOR2X1 U658 (.IN1(round_key[72]), .IN2(block[72]), .Q(n645));
   AO221X1 U659 (.IN1(n777), .IN2(n650), .IN3(n453), .IN4(new_block[71]), .IN5(n651), .Q(
          n1172));
   AO222X1 U660 (.IN1(n770), .IN2(new_sboxw[7]), .IN3(n1016), .IN4(n652), .IN5(n1259), .
          IN6(n653), .Q(n651));
   XOR3X1 U661 (.IN1(n654), .IN2(n237), .IN3(n655), .Q(n653));
   XOR2X1 U663 (.IN1(new_block[55]), .IN2(new_block[15]), .Q(n654));
   XOR2X1 U664 (.IN1(round_key[71]), .IN2(new_block[103]), .Q(n652));
   XOR2X1 U665 (.IN1(round_key[71]), .IN2(block[71]), .Q(n650));
   AO221X1 U666 (.IN1(n827), .IN2(n656), .IN3(n453), .IN4(new_block[70]), .IN5(n657), .Q(
          n1173));
   AO222X1 U667 (.IN1(n770), .IN2(new_sboxw[6]), .IN3(n1023), .IN4(n658), .IN5(n1258), .
          IN6(n659), .Q(n657));
   XOR3X1 U668 (.IN1(n660), .IN2(n238), .IN3(n661), .Q(n659));
   XOR3X1 U669 (.IN1(round_key[70]), .IN2(new_block[94]), .IN3(n206), .Q(n661));
   XOR2X1 U670 (.IN1(new_block[54]), .IN2(new_block[14]), .Q(n660));
   XOR2X1 U671 (.IN1(round_key[70]), .IN2(new_block[102]), .Q(n658));
   XOR2X1 U672 (.IN1(round_key[70]), .IN2(block[70]), .Q(n656));
   AO221X1 U673 (.IN1(n790), .IN2(n662), .IN3(n453), .IN4(new_block[69]), .IN5(n663), .Q(
          n1174));
   AO222X1 U674 (.IN1(n770), .IN2(new_sboxw[5]), .IN3(n986), .IN4(n664), .IN5(n1259), .IN6(
          n665), .Q(n663));
   XOR3X1 U675 (.IN1(n666), .IN2(n239), .IN3(n667), .Q(n665));
   XOR3X1 U676 (.IN1(round_key[69]), .IN2(new_block[93]), .IN3(n207), .Q(n667));
   XOR2X1 U677 (.IN1(new_block[53]), .IN2(new_block[13]), .Q(n666));
   XOR2X1 U678 (.IN1(round_key[69]), .IN2(new_block[101]), .Q(n664));
   XOR2X1 U679 (.IN1(round_key[69]), .IN2(block[69]), .Q(n662));
   AO221X1 U680 (.IN1(n966), .IN2(n668), .IN3(n453), .IN4(new_block[68]), .IN5(n669), .Q(
          n1175));
   AO222X1 U681 (.IN1(n701), .IN2(new_sboxw[4]), .IN3(n986), .IN4(n670), .IN5(n1261), .IN6(
          n671), .Q(n669));
   XNOR3X1 U683 (.IN1(n524), .IN2(new_block[12]), .IN3(n624), .Q(n673));
   XOR2X1 U684 (.IN1(n240), .IN2(new_block[103]), .Q(n624));
   XOR2X1 U685 (.IN1(new_block[91]), .IN2(new_block[95]), .Q(n524));
   XOR2X1 U687 (.IN1(round_key[68]), .IN2(new_block[100]), .Q(n670));
   XOR2X1 U688 (.IN1(round_key[68]), .IN2(block[68]), .Q(n668));
   AO221X1 U689 (.IN1(n790), .IN2(n674), .IN3(n453), .IN4(new_block[67]), .IN5(n675), .Q(
          n1176));
   AO222X1 U690 (.IN1(n770), .IN2(new_sboxw[3]), .IN3(n1036), .IN4(n676), .IN5(n1259), .
          IN6(n677), .Q(n675));
   XOR3X1 U692 (.IN1(n531), .IN2(n167), .IN3(n631), .Q(n679));
   XOR2X1 U693 (.IN1(n241), .IN2(new_block[103]), .Q(n631));
   XOR2X1 U694 (.IN1(new_block[90]), .IN2(new_block[95]), .Q(n531));
   XOR2X1 U696 (.IN1(round_key[67]), .IN2(new_block[99]), .Q(n676));
   XOR2X1 U697 (.IN1(round_key[67]), .IN2(block[67]), .Q(n674));
   AO221X1 U698 (.IN1(n820), .IN2(n680), .IN3(n453), .IN4(new_block[66]), .IN5(n681), .Q(
          n1177));
   AO222X1 U699 (.IN1(n701), .IN2(new_sboxw[2]), .IN3(n1036), .IN4(n682), .IN5(n1259), .
          IN6(n683), .Q(n681));
   XOR3X1 U700 (.IN1(n684), .IN2(n168), .IN3(n685), .Q(n683));
   XNOR3X1 U701 (.IN1(round_key[66]), .IN2(new_block[97]), .IN3(new_block[90]), .Q(n685)
          );
   XOR2X1 U702 (.IN1(new_block[89]), .IN2(new_block[50]), .Q(n684));
   XOR2X1 U703 (.IN1(round_key[66]), .IN2(new_block[98]), .Q(n682));
   XOR2X1 U704 (.IN1(round_key[66]), .IN2(block[66]), .Q(n680));
   AO221X1 U705 (.IN1(n870), .IN2(n686), .IN3(n453), .IN4(new_block[65]), .IN5(n687), .Q(
          n1178));
   AO222X1 U706 (.IN1(n770), .IN2(new_sboxw[1]), .IN3(n1023), .IN4(n688), .IN5(n1260), .
          IN6(n689), .Q(n687));
   XOR3X1 U708 (.IN1(n543), .IN2(n191), .IN3(n644), .Q(n691));
   XOR2X1 U709 (.IN1(new_block[96]), .IN2(n236), .Q(n644));
   XOR2X1 U711 (.IN1(round_key[65]), .IN2(new_block[97]), .Q(n688));
   XOR2X1 U712 (.IN1(round_key[65]), .IN2(block[65]), .Q(n686));
   AO221X1 U713 (.IN1(n840), .IN2(n692), .IN3(n453), .IN4(new_block[64]), .IN5(n693), .Q(
          n1179));
   AO222X1 U714 (.IN1(new_sboxw[0]), .IN2(n701), .IN3(n1036), .IN4(n694), .IN5(n433), .IN6(
          n695), .Q(n693));
   XOR3X1 U715 (.IN1(n543), .IN2(n236), .IN3(n696), .Q(n695));
   XNOR3X1 U716 (.IN1(round_key[64]), .IN2(new_block[8]), .IN3(new_block[48]), .Q(n696));
   XOR2X1 U717 (.IN1(new_block[88]), .IN2(new_block[95]), .Q(n543));
   XOR2X1 U718 (.IN1(round_key[64]), .IN2(new_block[96]), .Q(n694));
   XOR2X1 U720 (.IN1(round_key[64]), .IN2(block[64]), .Q(n692));
   AO221X1 U721 (.IN1(n678), .IN2(new_sboxw[31]), .IN3(n622), .IN4(new_block[63]), .IN5(
          n702), .Q(n1180));
   AO22X1 U722 (.IN1(round_key[63]), .IN2(n703), .IN3(n704), .IN4(n1299), .Q(n702));
   AO222X1 U723 (.IN1(block[63]), .IN2(n840), .IN3(n1257), .IN4(n705), .IN5(n1254), .IN6(
          new_block[63]), .Q(n704));
   OAI222X1 U724 (.IN1(n705), .IN2(n316), .IN3(n317), .IN4(new_block[63]), .IN5(n876), .
          IN6(block[63]), .QN(n703));
   XOR3X1 U725 (.IN1(new_block[22]), .IN2(n228), .IN3(n706), .Q(n705));
   XOR3X1 U726 (.IN1(new_block[71]), .IN2(new_block[62]), .IN3(n159), .Q(n706));
   AO221X1 U727 (.IN1(n678), .IN2(new_sboxw[30]), .IN3(n629), .IN4(new_block[62]), .IN5(
          n707), .Q(n1181));
   AO22X1 U728 (.IN1(round_key[62]), .IN2(n708), .IN3(n709), .IN4(n1300), .Q(n707));
   AO222X1 U729 (.IN1(block[62]), .IN2(n840), .IN3(n1264), .IN4(n710), .IN5(n973), .IN6(
          new_block[62]), .Q(n709));
   OAI222X1 U730 (.IN1(n710), .IN2(n1262), .IN3(n1084), .IN4(new_block[62]), .IN5(n318), .
          IN6(block[62]), .QN(n708));
   XOR3X1 U731 (.IN1(new_block[21]), .IN2(n229), .IN3(n711), .Q(n710));
   XOR3X1 U732 (.IN1(new_block[70]), .IN2(new_block[61]), .IN3(n160), .Q(n711));
   AO221X1 U733 (.IN1(n678), .IN2(new_sboxw[29]), .IN3(n622), .IN4(new_block[61]), .IN5(
          n712), .Q(n1182));
   AO22X1 U734 (.IN1(round_key[61]), .IN2(n713), .IN3(n714), .IN4(n1301), .Q(n712));
   AO222X1 U735 (.IN1(block[61]), .IN2(n777), .IN3(n1255), .IN4(n715), .IN5(n986), .IN6(
          new_block[61]), .Q(n714));
   OAI222X1 U736 (.IN1(n715), .IN2(n1262), .IN3(n1072), .IN4(new_block[61]), .IN5(n888), .
          IN6(block[61]), .QN(n713));
   XOR3X1 U737 (.IN1(new_block[20]), .IN2(n230), .IN3(n716), .Q(n715));
   XOR3X1 U738 (.IN1(new_block[69]), .IN2(new_block[60]), .IN3(n161), .Q(n716));
   AO221X1 U739 (.IN1(n678), .IN2(new_sboxw[28]), .IN3(n629), .IN4(new_block[60]), .IN5(
          n717), .Q(n1183));
   AO22X1 U740 (.IN1(round_key[60]), .IN2(n718), .IN3(n719), .IN4(n1302), .Q(n717));
   AO222X1 U741 (.IN1(block[60]), .IN2(n870), .IN3(n1255), .IN4(n720), .IN5(n1036), .IN6(
          new_block[60]), .Q(n719));
   OAI222X1 U742 (.IN1(n720), .IN2(n1263), .IN3(n1084), .IN4(new_block[60]), .IN5(n876), .
          IN6(block[60]), .QN(n718));
   XNOR3X1 U743 (.IN1(n721), .IN2(n722), .IN3(n723), .Q(n720));
   XOR3X1 U744 (.IN1(new_block[68]), .IN2(new_block[20]), .IN3(n231), .Q(n723));
   AO221X1 U745 (.IN1(n678), .IN2(new_sboxw[27]), .IN3(n622), .IN4(new_block[59]), .IN5(
          n724), .Q(n1184));
   AO22X1 U746 (.IN1(round_key[59]), .IN2(n725), .IN3(n726), .IN4(n1303), .Q(n724));
   AO222X1 U747 (.IN1(block[59]), .IN2(n840), .IN3(n1255), .IN4(n727), .IN5(n986), .IN6(
          new_block[59]), .Q(n726));
   OAI222X1 U748 (.IN1(n727), .IN2(n1262), .IN3(n1072), .IN4(new_block[59]), .IN5(n876), .
          IN6(block[59]), .QN(n725));
   XNOR3X1 U749 (.IN1(n728), .IN2(n729), .IN3(n730), .Q(n727));
   XOR3X1 U750 (.IN1(new_block[67]), .IN2(new_block[19]), .IN3(n232), .Q(n730));
   AO221X1 U751 (.IN1(n678), .IN2(new_sboxw[26]), .IN3(n629), .IN4(new_block[58]), .IN5(
          n731), .Q(n1185));
   AO22X1 U752 (.IN1(round_key[58]), .IN2(n732), .IN3(n733), .IN4(n1304), .Q(n731));
   AO222X1 U753 (.IN1(block[58]), .IN2(n840), .IN3(n1255), .IN4(n734), .IN5(n1066), .IN6(
          new_block[58]), .Q(n733));
   OAI222X1 U754 (.IN1(n734), .IN2(n1262), .IN3(n317), .IN4(new_block[58]), .IN5(n318), .
          IN6(block[58]), .QN(n732));
   XOR3X1 U755 (.IN1(new_block[17]), .IN2(n233), .IN3(n735), .Q(n734));
   XOR3X1 U756 (.IN1(new_block[66]), .IN2(new_block[57]), .IN3(n164), .Q(n735));
   AO221X1 U757 (.IN1(n678), .IN2(new_sboxw[25]), .IN3(n622), .IN4(new_block[57]), .IN5(
          n736), .Q(n1186));
   AO22X1 U758 (.IN1(round_key[57]), .IN2(n737), .IN3(n738), .IN4(n1305), .Q(n736));
   AO222X1 U759 (.IN1(block[57]), .IN2(n820), .IN3(n1258), .IN4(n739), .IN5(n1016), .IN6(
          new_block[57]), .Q(n738));
   OAI222X1 U760 (.IN1(n739), .IN2(n1263), .IN3(n1072), .IN4(new_block[57]), .IN5(n318), .
          IN6(block[57]), .QN(n737));
   XNOR3X1 U761 (.IN1(n740), .IN2(n741), .IN3(n742), .Q(n739));
   XOR3X1 U762 (.IN1(new_block[65]), .IN2(new_block[17]), .IN3(n234), .Q(n742));
   AO221X1 U763 (.IN1(n678), .IN2(new_sboxw[24]), .IN3(n629), .IN4(new_block[56]), .IN5(
          n743), .Q(n1187));
   AO22X1 U764 (.IN1(round_key[56]), .IN2(n744), .IN3(n745), .IN4(n1306), .Q(n743));
   AO222X1 U765 (.IN1(block[56]), .IN2(n390), .IN3(n1257), .IN4(n746), .IN5(n1113), .IN6(
          new_block[56]), .Q(n745));
   OAI222X1 U766 (.IN1(n746), .IN2(n1263), .IN3(n1084), .IN4(new_block[56]), .IN5(n318), .
          IN6(block[56]), .QN(n744));
   XOR3X1 U767 (.IN1(new_block[64]), .IN2(n181), .IN3(n747), .Q(n746));
   XOR2X1 U768 (.IN1(n235), .IN2(n740), .Q(n747));
   AO221X1 U769 (.IN1(n390), .IN2(n748), .IN3(n629), .IN4(new_block[55]), .IN5(n749), .Q(
          n1188));
   AO222X1 U770 (.IN1(n678), .IN2(new_sboxw[23]), .IN3(n1016), .IN4(n750), .IN5(n1264), .
          IN6(n751), .Q(n749));
   XOR3X1 U771 (.IN1(n752), .IN2(n229), .IN3(n753), .Q(n751));
   XOR3X1 U772 (.IN1(round_key[55]), .IN2(new_block[71]), .IN3(n181), .Q(n753));
   XOR2X1 U773 (.IN1(new_block[22]), .IN2(new_block[111]), .Q(n752));
   XOR2X1 U774 (.IN1(round_key[55]), .IN2(new_block[23]), .Q(n750));
   XOR2X1 U775 (.IN1(round_key[55]), .IN2(block[55]), .Q(n748));
   AO221X1 U776 (.IN1(n870), .IN2(n754), .IN3(n629), .IN4(new_block[54]), .IN5(n755), .Q(
          n1189));
   AO222X1 U777 (.IN1(n678), .IN2(new_sboxw[22]), .IN3(n973), .IN4(n756), .IN5(n1260), .
          IN6(n757), .Q(n755));
   XOR3X1 U778 (.IN1(n758), .IN2(n230), .IN3(n759), .Q(n757));
   XOR3X1 U779 (.IN1(round_key[54]), .IN2(new_block[70]), .IN3(n182), .Q(n759));
   XOR2X1 U780 (.IN1(new_block[21]), .IN2(new_block[110]), .Q(n758));
   XOR2X1 U781 (.IN1(round_key[54]), .IN2(new_block[22]), .Q(n756));
   XOR2X1 U782 (.IN1(round_key[54]), .IN2(block[54]), .Q(n754));
   AO221X1 U783 (.IN1(n966), .IN2(n760), .IN3(n629), .IN4(new_block[53]), .IN5(n761), .Q(
          n1190));
   AO222X1 U784 (.IN1(n678), .IN2(new_sboxw[21]), .IN3(n1023), .IN4(n762), .IN5(n1256), .
          IN6(n763), .Q(n761));
   XOR3X1 U785 (.IN1(n764), .IN2(n231), .IN3(n765), .Q(n763));
   XOR3X1 U786 (.IN1(round_key[53]), .IN2(new_block[69]), .IN3(n183), .Q(n765));
   XOR2X1 U787 (.IN1(new_block[20]), .IN2(new_block[109]), .Q(n764));
   XOR2X1 U788 (.IN1(round_key[53]), .IN2(new_block[21]), .Q(n762));
   XOR2X1 U789 (.IN1(round_key[53]), .IN2(block[53]), .Q(n760));
   AO221X1 U790 (.IN1(n897), .IN2(n766), .IN3(n629), .IN4(new_block[52]), .IN5(n767), .Q(
          n1191));
   AO222X1 U791 (.IN1(n678), .IN2(new_sboxw[20]), .IN3(n1066), .IN4(n768), .IN5(n433), .
          IN6(n769), .Q(n767));
   XOR3X1 U793 (.IN1(n721), .IN2(new_block[108]), .IN3(n772), .Q(n771));
   XOR2X1 U794 (.IN1(new_block[19]), .IN2(new_block[23]), .Q(n721));
   XOR2X1 U796 (.IN1(round_key[52]), .IN2(new_block[20]), .Q(n768));
   XOR2X1 U797 (.IN1(round_key[52]), .IN2(block[52]), .Q(n766));
   AO221X1 U798 (.IN1(n870), .IN2(n773), .IN3(n629), .IN4(new_block[51]), .IN5(n774), .Q(
          n1192));
   AO222X1 U799 (.IN1(n678), .IN2(new_sboxw[19]), .IN3(n403), .IN4(n775), .IN5(n1260), .
          IN6(n776), .Q(n774));
   XOR3X1 U801 (.IN1(n728), .IN2(new_block[107]), .IN3(n779), .Q(n778));
   XOR2X1 U802 (.IN1(new_block[18]), .IN2(new_block[23]), .Q(n728));
   XOR2X1 U804 (.IN1(round_key[51]), .IN2(new_block[19]), .Q(n775));
   XOR2X1 U805 (.IN1(round_key[51]), .IN2(block[51]), .Q(n773));
   AO221X1 U806 (.IN1(n840), .IN2(n780), .IN3(n629), .IN4(new_block[50]), .IN5(n781), .Q(
          n1193));
   AO222X1 U807 (.IN1(n690), .IN2(new_sboxw[18]), .IN3(n1113), .IN4(n782), .IN5(n1259), .
          IN6(n783), .Q(n781));
   XOR3X1 U808 (.IN1(n784), .IN2(n234), .IN3(n785), .Q(n783));
   XOR3X1 U809 (.IN1(round_key[50]), .IN2(new_block[66]), .IN3(n184), .Q(n785));
   XOR2X1 U810 (.IN1(new_block[17]), .IN2(new_block[106]), .Q(n784));
   XOR2X1 U811 (.IN1(round_key[50]), .IN2(new_block[18]), .Q(n782));
   XOR2X1 U812 (.IN1(round_key[50]), .IN2(block[50]), .Q(n780));
   AO221X1 U813 (.IN1(n777), .IN2(n786), .IN3(n629), .IN4(new_block[49]), .IN5(n787), .Q(
          n1194));
   AO222X1 U814 (.IN1(n690), .IN2(new_sboxw[17]), .IN3(n986), .IN4(n788), .IN5(n1257), .
          IN6(n789), .Q(n787));
   XOR3X1 U816 (.IN1(n740), .IN2(new_block[105]), .IN3(n792), .Q(n791));
   XOR2X1 U817 (.IN1(new_block[16]), .IN2(new_block[23]), .Q(n740));
   XOR2X1 U819 (.IN1(round_key[49]), .IN2(new_block[17]), .Q(n788));
   XOR2X1 U820 (.IN1(round_key[49]), .IN2(block[49]), .Q(n786));
   AO221X1 U821 (.IN1(n820), .IN2(n793), .IN3(n629), .IN4(new_block[48]), .IN5(n794), .Q(
          n1195));
   AO222X1 U822 (.IN1(n690), .IN2(new_sboxw[16]), .IN3(n973), .IN4(n795), .IN5(n1258), .
          IN6(n796), .Q(n794));
   XOR3X1 U823 (.IN1(n792), .IN2(n159), .IN3(n797), .Q(n796));
   XNOR3X1 U824 (.IN1(round_key[48]), .IN2(new_block[64]), .IN3(new_block[56]), .Q(n797)
          );
   XOR2X1 U825 (.IN1(round_key[48]), .IN2(new_block[16]), .Q(n795));
   XOR2X1 U826 (.IN1(round_key[48]), .IN2(block[48]), .Q(n793));
   AO221X1 U827 (.IN1(n790), .IN2(n798), .IN3(n629), .IN4(new_block[47]), .IN5(n799), .Q(
          n1196));
   AO222X1 U828 (.IN1(n690), .IN2(new_sboxw[15]), .IN3(n1066), .IN4(n800), .IN5(n1256), .
          IN6(n801), .Q(n799));
   XOR3X1 U829 (.IN1(n802), .IN2(n229), .IN3(n803), .Q(n801));
   XOR2X1 U831 (.IN1(new_block[63]), .IN2(new_block[23]), .Q(n802));
   XOR2X1 U832 (.IN1(round_key[47]), .IN2(new_block[111]), .Q(n800));
   XOR2X1 U833 (.IN1(round_key[47]), .IN2(block[47]), .Q(n798));
   AO221X1 U834 (.IN1(n827), .IN2(n804), .IN3(n629), .IN4(new_block[46]), .IN5(n805), .Q(
          n1197));
   AO222X1 U835 (.IN1(n690), .IN2(new_sboxw[14]), .IN3(n1016), .IN4(n806), .IN5(n1258), .
          IN6(n807), .Q(n805));
   XOR3X1 U836 (.IN1(n808), .IN2(n230), .IN3(n809), .Q(n807));
   XOR3X1 U837 (.IN1(round_key[46]), .IN2(new_block[70]), .IN3(n213), .Q(n809));
   XOR2X1 U838 (.IN1(new_block[62]), .IN2(new_block[22]), .Q(n808));
   XOR2X1 U839 (.IN1(round_key[46]), .IN2(new_block[110]), .Q(n806));
   XOR2X1 U840 (.IN1(round_key[46]), .IN2(block[46]), .Q(n804));
   AO221X1 U841 (.IN1(n820), .IN2(n810), .IN3(n629), .IN4(new_block[45]), .IN5(n811), .Q(
          n1198));
   AO222X1 U842 (.IN1(n690), .IN2(new_sboxw[13]), .IN3(n1036), .IN4(n812), .IN5(n1259), .
          IN6(n813), .Q(n811));
   XOR3X1 U843 (.IN1(n814), .IN2(n231), .IN3(n815), .Q(n813));
   XOR3X1 U844 (.IN1(round_key[45]), .IN2(new_block[69]), .IN3(n214), .Q(n815));
   XOR2X1 U845 (.IN1(new_block[61]), .IN2(new_block[21]), .Q(n814));
   XOR2X1 U846 (.IN1(round_key[45]), .IN2(new_block[109]), .Q(n812));
   XOR2X1 U847 (.IN1(round_key[45]), .IN2(block[45]), .Q(n810));
   AO221X1 U848 (.IN1(n827), .IN2(n816), .IN3(n629), .IN4(new_block[44]), .IN5(n817), .Q(
          n1199));
   AO222X1 U849 (.IN1(n690), .IN2(new_sboxw[12]), .IN3(n973), .IN4(n818), .IN5(n433), .IN6(
          n819), .Q(n817));
   XOR3X1 U851 (.IN1(n772), .IN2(n162), .IN3(n822), .Q(n821));
   XOR2X1 U852 (.IN1(n232), .IN2(n228), .Q(n772));
   XOR2X1 U854 (.IN1(round_key[44]), .IN2(new_block[108]), .Q(n818));
   XOR2X1 U855 (.IN1(round_key[44]), .IN2(block[44]), .Q(n816));
   AO221X1 U856 (.IN1(n820), .IN2(n823), .IN3(n622), .IN4(new_block[43]), .IN5(n824), .Q(
          n1200));
   AO222X1 U857 (.IN1(n690), .IN2(new_sboxw[11]), .IN3(n1023), .IN4(n825), .IN5(n1260), .
          IN6(n826), .Q(n824));
   XOR3X1 U859 (.IN1(n779), .IN2(n163), .IN3(n829), .Q(n828));
   XOR2X1 U860 (.IN1(n233), .IN2(n228), .Q(n779));
   XOR2X1 U862 (.IN1(round_key[43]), .IN2(new_block[107]), .Q(n825));
   XOR2X1 U863 (.IN1(round_key[43]), .IN2(block[43]), .Q(n823));
   AO221X1 U864 (.IN1(n820), .IN2(n830), .IN3(n622), .IN4(new_block[42]), .IN5(n831), .Q(
          n1201));
   AO222X1 U865 (.IN1(n690), .IN2(new_sboxw[10]), .IN3(n1016), .IN4(n832), .IN5(n1260), .
          IN6(n833), .Q(n831));
   XOR3X1 U866 (.IN1(n834), .IN2(n234), .IN3(n835), .Q(n833));
   XOR3X1 U867 (.IN1(round_key[42]), .IN2(new_block[66]), .IN3(n217), .Q(n835));
   XOR2X1 U868 (.IN1(new_block[58]), .IN2(new_block[18]), .Q(n834));
   XOR2X1 U869 (.IN1(round_key[42]), .IN2(new_block[106]), .Q(n832));
   XOR2X1 U870 (.IN1(round_key[42]), .IN2(block[42]), .Q(n830));
   AO221X1 U871 (.IN1(n827), .IN2(n836), .IN3(n622), .IN4(new_block[41]), .IN5(n837), .Q(
          n1202));
   AO222X1 U872 (.IN1(n690), .IN2(new_sboxw[9]), .IN3(n1066), .IN4(n838), .IN5(n1257), .
          IN6(n839), .Q(n837));
   XOR3X1 U874 (.IN1(n792), .IN2(n165), .IN3(n842), .Q(n841));
   XOR2X1 U875 (.IN1(n235), .IN2(n228), .Q(n792));
   XOR2X1 U877 (.IN1(round_key[41]), .IN2(new_block[105]), .Q(n838));
   XOR2X1 U878 (.IN1(round_key[41]), .IN2(block[41]), .Q(n836));
   AO221X1 U879 (.IN1(n777), .IN2(n843), .IN3(n622), .IN4(new_block[40]), .IN5(n844), .Q(
          n1203));
   AO222X1 U880 (.IN1(n690), .IN2(new_sboxw[8]), .IN3(n1036), .IN4(n845), .IN5(n1258), .
          IN6(n846), .Q(n844));
   XOR3X1 U881 (.IN1(n842), .IN2(new_block[111]), .IN3(n847), .Q(n846));
   XNOR3X1 U882 (.IN1(round_key[40]), .IN2(new_block[56]), .IN3(new_block[16]), .Q(n847)
          );
   XOR2X1 U883 (.IN1(round_key[40]), .IN2(new_block[104]), .Q(n845));
   XOR2X1 U884 (.IN1(round_key[40]), .IN2(block[40]), .Q(n843));
   AO221X1 U885 (.IN1(n790), .IN2(n848), .IN3(n622), .IN4(new_block[39]), .IN5(n849), .Q(
          n1204));
   AO222X1 U886 (.IN1(n690), .IN2(new_sboxw[7]), .IN3(n973), .IN4(n850), .IN5(n1259), .IN6(
          n851), .Q(n849));
   XOR3X1 U887 (.IN1(n852), .IN2(n228), .IN3(n853), .Q(n851));
   XOR3X1 U888 (.IN1(round_key[39]), .IN2(new_block[70]), .IN3(n181), .Q(n853));
   XOR2X1 U889 (.IN1(new_block[62]), .IN2(new_block[23]), .Q(n852));
   XOR2X1 U890 (.IN1(round_key[39]), .IN2(new_block[71]), .Q(n850));
   XOR2X1 U891 (.IN1(round_key[39]), .IN2(block[39]), .Q(n848));
   AO221X1 U892 (.IN1(n790), .IN2(n854), .IN3(n622), .IN4(new_block[38]), .IN5(n855), .Q(
          n1205));
   AO222X1 U893 (.IN1(n690), .IN2(new_sboxw[6]), .IN3(n1023), .IN4(n856), .IN5(n1261), .
          IN6(n857), .Q(n855));
   XOR3X1 U894 (.IN1(n858), .IN2(n229), .IN3(n859), .Q(n857));
   XOR3X1 U895 (.IN1(round_key[38]), .IN2(new_block[69]), .IN3(n182), .Q(n859));
   XOR2X1 U896 (.IN1(new_block[61]), .IN2(new_block[22]), .Q(n858));
   XOR2X1 U897 (.IN1(round_key[38]), .IN2(new_block[70]), .Q(n856));
   XOR2X1 U898 (.IN1(round_key[38]), .IN2(block[38]), .Q(n854));
   AO221X1 U899 (.IN1(n777), .IN2(n860), .IN3(n622), .IN4(new_block[37]), .IN5(n861), .Q(
          n1206));
   AO222X1 U900 (.IN1(n690), .IN2(new_sboxw[5]), .IN3(n1254), .IN4(n862), .IN5(n1259), .
          IN6(n863), .Q(n861));
   XOR3X1 U901 (.IN1(n864), .IN2(n230), .IN3(n865), .Q(n863));
   XOR3X1 U902 (.IN1(round_key[37]), .IN2(new_block[68]), .IN3(n183), .Q(n865));
   XOR2X1 U903 (.IN1(new_block[60]), .IN2(new_block[21]), .Q(n864));
   XOR2X1 U904 (.IN1(round_key[37]), .IN2(new_block[69]), .Q(n862));
   XOR2X1 U905 (.IN1(round_key[37]), .IN2(block[37]), .Q(n860));
   AO221X1 U906 (.IN1(n390), .IN2(n866), .IN3(n622), .IN4(new_block[36]), .IN5(n867), .Q(
          n1207));
   AO222X1 U907 (.IN1(n678), .IN2(new_sboxw[4]), .IN3(n1254), .IN4(n868), .IN5(n1256), .
          IN6(n869), .Q(n867));
   XOR3X1 U909 (.IN1(n722), .IN2(n231), .IN3(n822), .Q(n871));
   XOR2X1 U910 (.IN1(n215), .IN2(new_block[71]), .Q(n822));
   XOR2X1 U911 (.IN1(new_block[59]), .IN2(new_block[63]), .Q(n722));
   XOR2X1 U913 (.IN1(round_key[36]), .IN2(new_block[68]), .Q(n868));
   XOR2X1 U914 (.IN1(round_key[36]), .IN2(block[36]), .Q(n866));
   AO221X1 U915 (.IN1(n790), .IN2(n872), .IN3(n622), .IN4(new_block[35]), .IN5(n873), .Q(
          n1208));
   AO222X1 U916 (.IN1(n678), .IN2(new_sboxw[3]), .IN3(n403), .IN4(n874), .IN5(n1260), .IN6(
          n875), .Q(n873));
   XOR3X1 U918 (.IN1(n729), .IN2(n232), .IN3(n829), .Q(n877));
   XOR2X1 U919 (.IN1(n216), .IN2(new_block[71]), .Q(n829));
   XOR2X1 U920 (.IN1(new_block[58]), .IN2(new_block[63]), .Q(n729));
   XOR2X1 U922 (.IN1(round_key[35]), .IN2(new_block[67]), .Q(n874));
   XOR2X1 U923 (.IN1(round_key[35]), .IN2(block[35]), .Q(n872));
   AO221X1 U924 (.IN1(n966), .IN2(n878), .IN3(n622), .IN4(new_block[34]), .IN5(n879), .Q(
          n1209));
   AO222X1 U925 (.IN1(n678), .IN2(new_sboxw[2]), .IN3(n1016), .IN4(n880), .IN5(n1257), .
          IN6(n881), .Q(n879));
   XOR3X1 U926 (.IN1(n882), .IN2(n233), .IN3(n883), .Q(n881));
   XOR3X1 U927 (.IN1(round_key[34]), .IN2(new_block[65]), .IN3(n184), .Q(n883));
   XOR2X1 U928 (.IN1(new_block[57]), .IN2(new_block[18]), .Q(n882));
   XOR2X1 U929 (.IN1(round_key[34]), .IN2(new_block[66]), .Q(n880));
   XOR2X1 U930 (.IN1(round_key[34]), .IN2(block[34]), .Q(n878));
   AO221X1 U931 (.IN1(n897), .IN2(n884), .IN3(n622), .IN4(new_block[33]), .IN5(n885), .Q(
          n1210));
   AO222X1 U932 (.IN1(n690), .IN2(new_sboxw[1]), .IN3(n1016), .IN4(n886), .IN5(n1261), .
          IN6(n887), .Q(n885));
   XOR3X1 U934 (.IN1(n741), .IN2(n234), .IN3(n842), .Q(n889));
   XNOR2X1 U935 (.IN1(new_block[64]), .IN2(new_block[71]), .Q(n842));
   XOR2X1 U937 (.IN1(round_key[33]), .IN2(new_block[65]), .Q(n886));
   XOR2X1 U938 (.IN1(round_key[33]), .IN2(block[33]), .Q(n884));
   AO221X1 U939 (.IN1(n777), .IN2(n890), .IN3(n622), .IN4(new_block[32]), .IN5(n891), .Q(
          n1211));
   AO222X1 U940 (.IN1(n690), .IN2(new_sboxw[0]), .IN3(n1113), .IN4(n892), .IN5(n1264), .
          IN6(n893), .Q(n891));
   XOR3X1 U941 (.IN1(n741), .IN2(n235), .IN3(n894), .Q(n893));
   XNOR3X1 U942 (.IN1(round_key[32]), .IN2(new_block[71]), .IN3(new_block[16]), .Q(n894)
          );
   XOR2X1 U943 (.IN1(new_block[56]), .IN2(new_block[63]), .Q(n741));
   XOR2X1 U944 (.IN1(round_key[32]), .IN2(new_block[64]), .Q(n892));
   XOR2X1 U946 (.IN1(round_key[32]), .IN2(block[32]), .Q(n890));
   AO221X1 U947 (.IN1(n642), .IN2(new_sboxw[31]), .IN3(n501), .IN4(new_block[31]), .IN5(
          n898), .Q(n1212));
   AO22X1 U948 (.IN1(round_key[31]), .IN2(n899), .IN3(n900), .IN4(n1307), .Q(n898));
   AO222X1 U949 (.IN1(block[31]), .IN2(n966), .IN3(n1256), .IN4(n901), .IN5(n1113), .IN6(
          new_block[31]), .Q(n900));
   OAI222X1 U950 (.IN1(n901), .IN2(n316), .IN3(n1084), .IN4(new_block[31]), .IN5(n318), .
          IN6(block[31]), .QN(n899));
   XOR3X1 U951 (.IN1(new_block[119]), .IN2(n223), .IN3(n902), .Q(n901));
   XOR3X1 U952 (.IN1(new_block[79]), .IN2(n197), .IN3(new_block[30]), .Q(n902));
   AO221X1 U953 (.IN1(n642), .IN2(new_sboxw[30]), .IN3(n503), .IN4(new_block[30]), .IN5(
          n903), .Q(n1213));
   AO22X1 U954 (.IN1(round_key[30]), .IN2(n904), .IN3(n905), .IN4(n1308), .Q(n903));
   AO222X1 U955 (.IN1(block[30]), .IN2(n897), .IN3(n433), .IN4(n906), .IN5(n1254), .IN6(
          new_block[30]), .Q(n905));
   OAI222X1 U956 (.IN1(n906), .IN2(n1262), .IN3(n317), .IN4(new_block[30]), .IN5(n318), .
          IN6(block[30]), .QN(n904));
   XOR3X1 U957 (.IN1(new_block[118]), .IN2(n224), .IN3(n907), .Q(n906));
   XOR3X1 U958 (.IN1(new_block[78]), .IN2(n198), .IN3(new_block[29]), .Q(n907));
   AO221X1 U959 (.IN1(n642), .IN2(new_sboxw[29]), .IN3(n501), .IN4(new_block[29]), .IN5(
          n908), .Q(n1214));
   AO22X1 U960 (.IN1(round_key[29]), .IN2(n909), .IN3(n910), .IN4(n1309), .Q(n908));
   AO222X1 U961 (.IN1(block[29]), .IN2(n390), .IN3(n1261), .IN4(n911), .IN5(n1066), .IN6(
          new_block[29]), .Q(n910));
   OAI222X1 U962 (.IN1(n911), .IN2(n1263), .IN3(n1084), .IN4(new_block[29]), .IN5(n318), .
          IN6(block[29]), .QN(n909));
   XOR3X1 U963 (.IN1(new_block[117]), .IN2(n225), .IN3(n912), .Q(n911));
   XOR3X1 U964 (.IN1(new_block[77]), .IN2(n199), .IN3(new_block[28]), .Q(n912));
   AO221X1 U965 (.IN1(n642), .IN2(new_sboxw[28]), .IN3(n503), .IN4(new_block[28]), .IN5(
          n913), .Q(n1215));
   AO22X1 U966 (.IN1(round_key[28]), .IN2(n914), .IN3(n915), .IN4(n1310), .Q(n913));
   AO222X1 U967 (.IN1(block[28]), .IN2(n966), .IN3(n1264), .IN4(n916), .IN5(n403), .IN6(
          new_block[28]), .Q(n915));
   OAI222X1 U968 (.IN1(n916), .IN2(n1263), .IN3(n1084), .IN4(new_block[28]), .IN5(n318), .
          IN6(block[28]), .QN(n914));
   XNOR3X1 U969 (.IN1(n917), .IN2(n918), .IN3(n919), .Q(n916));
   XOR3X1 U970 (.IN1(new_block[76]), .IN2(new_block[36]), .IN3(n225), .Q(n919));
   AO221X1 U971 (.IN1(n642), .IN2(new_sboxw[27]), .IN3(n501), .IN4(new_block[27]), .IN5(
          n920), .Q(n1216));
   AO22X1 U972 (.IN1(round_key[27]), .IN2(n921), .IN3(n922), .IN4(n1311), .Q(n920));
   AO222X1 U973 (.IN1(block[27]), .IN2(n870), .IN3(n433), .IN4(n923), .IN5(n986), .IN6(
          new_block[27]), .Q(n922));
   OAI222X1 U974 (.IN1(n923), .IN2(n316), .IN3(n1084), .IN4(new_block[27]), .IN5(n318), .
          IN6(block[27]), .QN(n921));
   XNOR3X1 U975 (.IN1(n924), .IN2(n925), .IN3(n926), .Q(n923));
   XOR3X1 U976 (.IN1(new_block[75]), .IN2(new_block[35]), .IN3(n226), .Q(n926));
   AO221X1 U977 (.IN1(n642), .IN2(new_sboxw[26]), .IN3(n503), .IN4(new_block[26]), .IN5(
          n927), .Q(n1217));
   AO22X1 U978 (.IN1(round_key[26]), .IN2(n928), .IN3(n929), .IN4(n1312), .Q(n927));
   AO222X1 U979 (.IN1(block[26]), .IN2(n827), .IN3(n1261), .IN4(n930), .IN5(n1113), .IN6(
          new_block[26]), .Q(n929));
   OAI222X1 U980 (.IN1(n930), .IN2(n1262), .IN3(n1072), .IN4(new_block[26]), .IN5(n318), .
          IN6(block[26]), .QN(n928));
   XOR3X1 U981 (.IN1(new_block[114]), .IN2(n227), .IN3(n931), .Q(n930));
   XOR3X1 U982 (.IN1(new_block[74]), .IN2(n202), .IN3(new_block[25]), .Q(n931));
   AO221X1 U983 (.IN1(n642), .IN2(new_sboxw[25]), .IN3(n501), .IN4(new_block[25]), .IN5(
          n932), .Q(n1218));
   AO22X1 U984 (.IN1(round_key[25]), .IN2(n933), .IN3(n934), .IN4(n1313), .Q(n932));
   AO222X1 U985 (.IN1(block[25]), .IN2(n870), .IN3(n1256), .IN4(n935), .IN5(n973), .IN6(
          new_block[25]), .Q(n934));
   OAI222X1 U986 (.IN1(n935), .IN2(n1262), .IN3(n317), .IN4(new_block[25]), .IN5(n888), .
          IN6(block[25]), .QN(n933));
   XNOR3X1 U987 (.IN1(n936), .IN2(n937), .IN3(n938), .Q(n935));
   XOR3X1 U988 (.IN1(new_block[73]), .IN2(new_block[33]), .IN3(n227), .Q(n938));
   AO221X1 U989 (.IN1(n642), .IN2(new_sboxw[24]), .IN3(n503), .IN4(new_block[24]), .IN5(
          n939), .Q(n1219));
   AO22X1 U990 (.IN1(round_key[24]), .IN2(n940), .IN3(n941), .IN4(n1314), .Q(n939));
   AO222X1 U991 (.IN1(block[24]), .IN2(n820), .IN3(n1258), .IN4(n942), .IN5(n986), .IN6(
          new_block[24]), .Q(n941));
   OAI222X1 U992 (.IN1(n942), .IN2(n1263), .IN3(n1072), .IN4(new_block[24]), .IN5(n318), .
          IN6(block[24]), .QN(n940));
   XOR3X1 U993 (.IN1(new_block[72]), .IN2(n204), .IN3(n943), .Q(n942));
   XNOR2X1 U994 (.IN1(new_block[31]), .IN2(n936), .Q(n943));
   AO221X1 U995 (.IN1(n897), .IN2(n944), .IN3(n503), .IN4(new_block[23]), .IN5(n945), .Q(
          n1220));
   AO222X1 U996 (.IN1(n642), .IN2(new_sboxw[23]), .IN3(n973), .IN4(n946), .IN5(n1257), .
          IN6(n947), .Q(n945));
   XOR3X1 U997 (.IN1(n948), .IN2(n223), .IN3(n949), .Q(n947));
   XNOR3X1 U998 (.IN1(round_key[23]), .IN2(new_block[79]), .IN3(new_block[78]), .Q(n949)
          );
   XOR2X1 U999 (.IN1(new_block[39]), .IN2(new_block[31]), .Q(n948));
   XOR2X1 U1000 (.IN1(round_key[23]), .IN2(new_block[119]), .Q(n946));
   XOR2X1 U1001 (.IN1(round_key[23]), .IN2(block[23]), .Q(n944));
   AO221X1 U1002 (.IN1(n966), .IN2(n950), .IN3(n503), .IN4(new_block[22]), .IN5(n951), .Q(
          n1221));
   AO222X1 U1003 (.IN1(n642), .IN2(new_sboxw[22]), .IN3(n1036), .IN4(n952), .IN5(n1264), .
          IN6(n953), .Q(n951));
   XOR3X1 U1004 (.IN1(n954), .IN2(n224), .IN3(n955), .Q(n953));
   XNOR3X1 U1005 (.IN1(round_key[22]), .IN2(new_block[78]), .IN3(new_block[77]), .Q(n955)
          );
   XOR2X1 U1006 (.IN1(new_block[38]), .IN2(new_block[30]), .Q(n954));
   XOR2X1 U1007 (.IN1(round_key[22]), .IN2(new_block[118]), .Q(n952));
   XOR2X1 U1008 (.IN1(round_key[22]), .IN2(block[22]), .Q(n950));
   AO221X1 U1009 (.IN1(n840), .IN2(n956), .IN3(n503), .IN4(new_block[21]), .IN5(n957), .Q(
          n1222));
   AO222X1 U1010 (.IN1(n642), .IN2(new_sboxw[21]), .IN3(n1016), .IN4(n958), .IN5(n1258), .
          IN6(n959), .Q(n957));
   XOR3X1 U1011 (.IN1(n960), .IN2(n225), .IN3(n961), .Q(n959));
   XOR3X1 U1012 (.IN1(round_key[21]), .IN2(new_block[77]), .IN3(n208), .Q(n961));
   XOR2X1 U1013 (.IN1(new_block[37]), .IN2(new_block[29]), .Q(n960));
   XOR2X1 U1014 (.IN1(round_key[21]), .IN2(new_block[117]), .Q(n958));
   XOR2X1 U1015 (.IN1(round_key[21]), .IN2(block[21]), .Q(n956));
   AO221X1 U1016 (.IN1(n870), .IN2(n962), .IN3(n503), .IN4(new_block[20]), .IN5(n963), .Q(
          n1223));
   AO222X1 U1017 (.IN1(n642), .IN2(new_sboxw[20]), .IN3(n986), .IN4(n964), .IN5(n1259), .
          IN6(n965), .Q(n963));
   XOR3X1 U1019 (.IN1(n917), .IN2(new_block[28]), .IN3(n968), .Q(n967));
   XOR2X1 U1020 (.IN1(new_block[115]), .IN2(new_block[119]), .Q(n917));
   XOR2X1 U1022 (.IN1(round_key[20]), .IN2(new_block[116]), .Q(n964));
   XOR2X1 U1023 (.IN1(round_key[20]), .IN2(block[20]), .Q(n962));
   AO221X1 U1024 (.IN1(n390), .IN2(n969), .IN3(n503), .IN4(new_block[19]), .IN5(n970), .Q(
          n1224));
   AO222X1 U1025 (.IN1(n642), .IN2(new_sboxw[19]), .IN3(n973), .IN4(n971), .IN5(n1258), .
          IN6(n972), .Q(n970));
   XOR3X1 U1027 (.IN1(n924), .IN2(new_block[27]), .IN3(n975), .Q(n974));
   XOR2X1 U1028 (.IN1(new_block[114]), .IN2(new_block[119]), .Q(n924));
   XOR2X1 U1030 (.IN1(round_key[19]), .IN2(new_block[115]), .Q(n971));
   XOR2X1 U1031 (.IN1(round_key[19]), .IN2(block[19]), .Q(n969));
   AO221X1 U1032 (.IN1(n790), .IN2(n976), .IN3(n503), .IN4(new_block[18]), .IN5(n977), .Q(
          n1225));
   AO222X1 U1033 (.IN1(n642), .IN2(new_sboxw[18]), .IN3(n1113), .IN4(n978), .IN5(n1261), .
          IN6(n979), .Q(n977));
   XOR3X1 U1034 (.IN1(n980), .IN2(n227), .IN3(n981), .Q(n979));
   XOR3X1 U1035 (.IN1(round_key[18]), .IN2(new_block[74]), .IN3(n210), .Q(n981));
   XOR2X1 U1036 (.IN1(new_block[34]), .IN2(new_block[26]), .Q(n980));
   XOR2X1 U1037 (.IN1(round_key[18]), .IN2(new_block[114]), .Q(n978));
   XOR2X1 U1038 (.IN1(round_key[18]), .IN2(block[18]), .Q(n976));
   AO221X1 U1039 (.IN1(n777), .IN2(n982), .IN3(n503), .IN4(new_block[17]), .IN5(n983), .Q(
          n1226));
   AO222X1 U1040 (.IN1(n672), .IN2(new_sboxw[17]), .IN3(n1254), .IN4(n984), .IN5(n1264), .
          IN6(n985), .Q(n983));
   XOR3X1 U1042 (.IN1(n936), .IN2(new_block[25]), .IN3(n988), .Q(n987));
   XOR2X1 U1043 (.IN1(new_block[112]), .IN2(new_block[119]), .Q(n936));
   XOR2X1 U1045 (.IN1(round_key[17]), .IN2(new_block[113]), .Q(n984));
   XOR2X1 U1046 (.IN1(round_key[17]), .IN2(block[17]), .Q(n982));
   AO221X1 U1047 (.IN1(n827), .IN2(n989), .IN3(n503), .IN4(new_block[16]), .IN5(n990), .Q(
          n1227));
   AO222X1 U1048 (.IN1(n642), .IN2(new_sboxw[16]), .IN3(n403), .IN4(n991), .IN5(n1256), .
          IN6(n992), .Q(n990));
   XNOR3X1 U1049 (.IN1(n988), .IN2(new_block[119]), .IN3(n993), .Q(n992));
   XOR3X1 U1050 (.IN1(round_key[16]), .IN2(n204), .IN3(new_block[24]), .Q(n993));
   XOR2X1 U1051 (.IN1(round_key[16]), .IN2(new_block[112]), .Q(n991));
   XOR2X1 U1052 (.IN1(round_key[16]), .IN2(block[16]), .Q(n989));
   AO221X1 U1053 (.IN1(n827), .IN2(n994), .IN3(n503), .IN4(new_block[15]), .IN5(n995), .Q(
          n1228));
   AO222X1 U1054 (.IN1(n672), .IN2(new_sboxw[15]), .IN3(n1023), .IN4(n996), .IN5(n1259), .
          IN6(n997), .Q(n995));
   XNOR3X1 U1055 (.IN1(n998), .IN2(new_block[119]), .IN3(n999), .Q(n997));
   XOR3X1 U1056 (.IN1(round_key[15]), .IN2(new_block[78]), .IN3(n197), .Q(n999));
   XOR2X1 U1057 (.IN1(new_block[38]), .IN2(new_block[31]), .Q(n998));
   XOR2X1 U1058 (.IN1(round_key[15]), .IN2(new_block[79]), .Q(n996));
   XOR2X1 U1059 (.IN1(round_key[15]), .IN2(block[15]), .Q(n994));
   AO221X1 U1060 (.IN1(n820), .IN2(n1000), .IN3(n503), .IN4(new_block[14]), .IN5(n1001), .
          Q(n1229));
   AO222X1 U1061 (.IN1(n672), .IN2(new_sboxw[14]), .IN3(n1023), .IN4(n1002), .IN5(n1255), .
          IN6(n1003), .Q(n1001));
   XOR3X1 U1062 (.IN1(n1004), .IN2(n223), .IN3(n1005), .Q(n1003));
   XOR3X1 U1063 (.IN1(round_key[14]), .IN2(new_block[77]), .IN3(n198), .Q(n1005));
   XOR2X1 U1064 (.IN1(new_block[37]), .IN2(new_block[30]), .Q(n1004));
   XOR2X1 U1065 (.IN1(round_key[14]), .IN2(new_block[78]), .Q(n1002));
   XOR2X1 U1066 (.IN1(round_key[14]), .IN2(block[14]), .Q(n1000));
   AO221X1 U1067 (.IN1(n870), .IN2(n1006), .IN3(n503), .IN4(new_block[13]), .IN5(n1007), .
          Q(n1230));
   AO222X1 U1068 (.IN1(n672), .IN2(new_sboxw[13]), .IN3(n403), .IN4(n1008), .IN5(n1261), .
          IN6(n1009), .Q(n1007));
   XOR3X1 U1069 (.IN1(n1010), .IN2(n224), .IN3(n1011), .Q(n1009));
   XOR3X1 U1070 (.IN1(round_key[13]), .IN2(new_block[76]), .IN3(n199), .Q(n1011));
   XOR2X1 U1071 (.IN1(new_block[36]), .IN2(new_block[29]), .Q(n1010));
   XOR2X1 U1072 (.IN1(round_key[13]), .IN2(new_block[77]), .Q(n1008));
   XOR2X1 U1073 (.IN1(round_key[13]), .IN2(block[13]), .Q(n1006));
   AO221X1 U1074 (.IN1(n840), .IN2(n1012), .IN3(n503), .IN4(new_block[12]), .IN5(n1013), .
          Q(n1231));
   AO222X1 U1075 (.IN1(n672), .IN2(new_sboxw[12]), .IN3(n1254), .IN4(n1014), .IN5(n1259), .
          IN6(n1015), .Q(n1013));
   XOR3X1 U1077 (.IN1(n968), .IN2(n225), .IN3(n1018), .Q(n1017));
   XNOR2X1 U1078 (.IN1(n209), .IN2(new_block[79]), .Q(n968));
   XOR2X1 U1080 (.IN1(round_key[12]), .IN2(new_block[76]), .Q(n1014));
   XOR2X1 U1081 (.IN1(round_key[12]), .IN2(block[12]), .Q(n1012));
   AO221X1 U1082 (.IN1(n870), .IN2(n1019), .IN3(n501), .IN4(new_block[11]), .IN5(n1020), .
          Q(n1232));
   AO222X1 U1083 (.IN1(n672), .IN2(new_sboxw[11]), .IN3(n1254), .IN4(n1021), .IN5(n1256), .
          IN6(n1022), .Q(n1020));
   XOR3X1 U1085 (.IN1(n975), .IN2(n226), .IN3(n1025), .Q(n1024));
   XOR2X1 U1086 (.IN1(new_block[74]), .IN2(new_block[79]), .Q(n975));
   XOR2X1 U1088 (.IN1(round_key[11]), .IN2(new_block[75]), .Q(n1021));
   XOR2X1 U1089 (.IN1(round_key[11]), .IN2(block[11]), .Q(n1019));
   AO221X1 U1090 (.IN1(n897), .IN2(n1026), .IN3(n501), .IN4(new_block[10]), .IN5(n1027), .
          Q(n1233));
   AO222X1 U1091 (.IN1(n672), .IN2(new_sboxw[10]), .IN3(n1254), .IN4(n1028), .IN5(n433), .
          IN6(n1029), .Q(n1027));
   XNOR3X1 U1092 (.IN1(n1030), .IN2(new_block[114]), .IN3(n1031), .Q(n1029));
   XOR3X1 U1093 (.IN1(round_key[10]), .IN2(new_block[73]), .IN3(n202), .Q(n1031));
   XOR2X1 U1094 (.IN1(new_block[33]), .IN2(new_block[26]), .Q(n1030));
   XOR2X1 U1095 (.IN1(round_key[10]), .IN2(new_block[74]), .Q(n1028));
   XOR2X1 U1096 (.IN1(round_key[10]), .IN2(block[10]), .Q(n1026));
   AO221X1 U1097 (.IN1(n966), .IN2(n1032), .IN3(n501), .IN4(new_block[9]), .IN5(n1033), .Q(
          n1234));
   AO222X1 U1098 (.IN1(n672), .IN2(new_sboxw[9]), .IN3(n1113), .IN4(n1034), .IN5(n1260), .
          IN6(n1035), .Q(n1033));
   XOR3X1 U1100 (.IN1(n988), .IN2(n227), .IN3(n1038), .Q(n1037));
   XNOR2X1 U1101 (.IN1(n211), .IN2(new_block[79]), .Q(n988));
   XOR2X1 U1103 (.IN1(round_key[9]), .IN2(new_block[73]), .Q(n1034));
   XOR2X1 U1104 (.IN1(round_key[9]), .IN2(block[9]), .Q(n1032));
   AO221X1 U1105 (.IN1(n390), .IN2(n1039), .IN3(n501), .IN4(new_block[8]), .IN5(n1040), .Q(
          n1235));
   AO222X1 U1106 (.IN1(n642), .IN2(new_sboxw[8]), .IN3(n986), .IN4(n1041), .IN5(n1257), .
          IN6(n1042), .Q(n1040));
   XOR3X1 U1107 (.IN1(n1038), .IN2(new_block[112]), .IN3(n1043), .Q(n1042));
   XNOR3X1 U1108 (.IN1(round_key[8]), .IN2(new_block[79]), .IN3(new_block[24]), .Q(n1043)
          );
   XOR2X1 U1109 (.IN1(round_key[8]), .IN2(new_block[72]), .Q(n1041));
   XOR2X1 U1110 (.IN1(round_key[8]), .IN2(block[8]), .Q(n1039));
   AO221X1 U1111 (.IN1(n897), .IN2(n1044), .IN3(n501), .IN4(new_block[7]), .IN5(n1045), .Q(
          n1236));
   AO222X1 U1112 (.IN1(n672), .IN2(new_sboxw[7]), .IN3(n1113), .IN4(n1046), .IN5(n1255), .
          IN6(n1047), .Q(n1045));
   XNOR3X1 U1113 (.IN1(n1048), .IN2(new_block[119]), .IN3(n1049), .Q(n1047));
   XOR3X1 U1114 (.IN1(round_key[7]), .IN2(new_block[79]), .IN3(n198), .Q(n1049));
   XOR2X1 U1115 (.IN1(new_block[31]), .IN2(new_block[30]), .Q(n1048));
   XOR2X1 U1116 (.IN1(round_key[7]), .IN2(new_block[39]), .Q(n1046));
   XOR2X1 U1117 (.IN1(round_key[7]), .IN2(block[7]), .Q(n1044));
   AO221X1 U1118 (.IN1(n966), .IN2(n1050), .IN3(n501), .IN4(new_block[6]), .IN5(n1051), .Q(
          n1237));
   AO222X1 U1119 (.IN1(n672), .IN2(new_sboxw[6]), .IN3(n1113), .IN4(n1052), .IN5(n1255), .
          IN6(n1053), .Q(n1051));
   XOR3X1 U1120 (.IN1(n1054), .IN2(n223), .IN3(n1055), .Q(n1053));
   XOR3X1 U1121 (.IN1(round_key[6]), .IN2(new_block[78]), .IN3(n199), .Q(n1055));
   XOR2X1 U1122 (.IN1(new_block[30]), .IN2(new_block[29]), .Q(n1054));
   XOR2X1 U1123 (.IN1(round_key[6]), .IN2(new_block[38]), .Q(n1052));
   XOR2X1 U1124 (.IN1(round_key[6]), .IN2(block[6]), .Q(n1050));
   AO221X1 U1125 (.IN1(n390), .IN2(n1056), .IN3(n501), .IN4(new_block[5]), .IN5(n1057), .Q(
          n1238));
   AO222X1 U1126 (.IN1(n672), .IN2(new_sboxw[5]), .IN3(n1066), .IN4(n1058), .IN5(n1256), .
          IN6(n1059), .Q(n1057));
   XOR3X1 U1127 (.IN1(n1060), .IN2(n224), .IN3(n1061), .Q(n1059));
   XOR3X1 U1128 (.IN1(round_key[5]), .IN2(new_block[77]), .IN3(n200), .Q(n1061));
   XOR2X1 U1129 (.IN1(new_block[29]), .IN2(new_block[28]), .Q(n1060));
   XOR2X1 U1130 (.IN1(round_key[5]), .IN2(new_block[37]), .Q(n1058));
   XOR2X1 U1131 (.IN1(round_key[5]), .IN2(block[5]), .Q(n1056));
   AO221X1 U1132 (.IN1(n966), .IN2(n1062), .IN3(n501), .IN4(new_block[4]), .IN5(n1063), .Q(
          n1239));
   AO222X1 U1133 (.IN1(n672), .IN2(new_sboxw[4]), .IN3(n1254), .IN4(n1064), .IN5(n433), .
          IN6(n1065), .Q(n1063));
   XOR3X1 U1135 (.IN1(n918), .IN2(n225), .IN3(n1018), .Q(n1067));
   XOR2X1 U1136 (.IN1(n201), .IN2(new_block[39]), .Q(n1018));
   XOR2X1 U1137 (.IN1(new_block[27]), .IN2(new_block[31]), .Q(n918));
   XOR2X1 U1139 (.IN1(round_key[4]), .IN2(new_block[36]), .Q(n1064));
   XOR2X1 U1140 (.IN1(round_key[4]), .IN2(block[4]), .Q(n1062));
   AO221X1 U1141 (.IN1(n827), .IN2(n1068), .IN3(n501), .IN4(new_block[3]), .IN5(n1069), .Q(
          n1240));
   AO222X1 U1142 (.IN1(n672), .IN2(new_sboxw[3]), .IN3(n1113), .IN4(n1070), .IN5(n1255), .
          IN6(n1071), .Q(n1069));
   XOR3X1 U1144 (.IN1(n925), .IN2(n226), .IN3(n1025), .Q(n1073));
   XOR2X1 U1145 (.IN1(n202), .IN2(new_block[39]), .Q(n1025));
   XOR2X1 U1146 (.IN1(new_block[26]), .IN2(new_block[31]), .Q(n925));
   XOR2X1 U1148 (.IN1(round_key[3]), .IN2(new_block[35]), .Q(n1070));
   XOR2X1 U1149 (.IN1(round_key[3]), .IN2(block[3]), .Q(n1068));
   AO221X1 U1150 (.IN1(n390), .IN2(n1074), .IN3(n501), .IN4(new_block[2]), .IN5(n1075), .Q(
          n1241));
   AO222X1 U1151 (.IN1(n672), .IN2(new_sboxw[2]), .IN3(n986), .IN4(n1076), .IN5(n1258), .
          IN6(n1077), .Q(n1075));
   XNOR3X1 U1152 (.IN1(n1078), .IN2(new_block[114]), .IN3(n1079), .Q(n1077));
   XOR3X1 U1153 (.IN1(round_key[2]), .IN2(new_block[74]), .IN3(n203), .Q(n1079));
   XOR2X1 U1154 (.IN1(new_block[26]), .IN2(new_block[25]), .Q(n1078));
   XOR2X1 U1155 (.IN1(round_key[2]), .IN2(new_block[34]), .Q(n1076));
   XOR2X1 U1156 (.IN1(round_key[2]), .IN2(block[2]), .Q(n1074));
   AO221X1 U1157 (.IN1(n390), .IN2(n1080), .IN3(n501), .IN4(new_block[1]), .IN5(n1081), .Q(
          n1242));
   AO222X1 U1158 (.IN1(n672), .IN2(new_sboxw[1]), .IN3(n1016), .IN4(n1082), .IN5(n1257), .
          IN6(n1083), .Q(n1081));
   XOR3X1 U1160 (.IN1(n937), .IN2(n227), .IN3(n1038), .Q(n1085));
   XOR2X1 U1161 (.IN1(new_block[32]), .IN2(n197), .Q(n1038));
   XOR2X1 U1163 (.IN1(round_key[1]), .IN2(new_block[33]), .Q(n1082));
   XOR2X1 U1164 (.IN1(round_key[1]), .IN2(block[1]), .Q(n1080));
   AO221X1 U1165 (.IN1(n827), .IN2(n1086), .IN3(n501), .IN4(new_block[0]), .IN5(n1087), .Q(
          n1243));
   AO222X1 U1166 (.IN1(n672), .IN2(new_sboxw[0]), .IN3(n1016), .IN4(n1088), .IN5(n433), .
          IN6(n1089), .Q(n1087));
   XNOR3X1 U1167 (.IN1(n937), .IN2(new_block[112]), .IN3(n1090), .Q(n1089));
   XOR3X1 U1168 (.IN1(round_key[0]), .IN2(new_block[72]), .IN3(n197), .Q(n1090));
   XOR2X1 U1169 (.IN1(new_block[24]), .IN2(new_block[31]), .Q(n937));
   XOR2X1 U1170 (.IN1(round_key[0]), .IN2(new_block[32]), .Q(n1088));
   XOR2X1 U1172 (.IN1(round_key[0]), .IN2(block[0]), .Q(n1086));
   AO221X1 U1173 (.IN1(n840), .IN2(n1093), .IN3(n579), .IN4(new_block[96]), .IN5(n1094), .
          Q(n1244));
   AO222X1 U1174 (.IN1(new_sboxw[0]), .IN2(n1266), .IN3(n973), .IN4(n1095), .IN5(n1261), .
          IN6(n1096), .Q(n1094));
   XOR3X1 U1175 (.IN1(n354), .IN2(n196), .IN3(n1097), .Q(n1096));
   XOR3X1 U1176 (.IN1(round_key[96]), .IN2(new_block[80]), .IN3(n169), .Q(n1097));
   XOR2X1 U1177 (.IN1(new_block[120]), .IN2(new_block[127]), .Q(n354));
   XOR2X1 U1178 (.IN1(round_key[96]), .IN2(new_block[0]), .Q(n1095));
   AND3X1 U1181 (.IN1(n318), .IN2(n317), .IN3(n316), .Q(n699));
   XOR2X1 U1182 (.IN1(round_key[96]), .IN2(block[96]), .Q(n1093));
   AO21X1 U1183 (.IN1(n1101), .IN2(n1102), .IN3(n1103), .Q(n1100));
   AO21X1 U1184 (.IN1(ready), .IN2(n1104), .IN3(n1036), .Q(n1245));
   OAI21X1 U1185 (.IN1(n1105), .IN2(n175), .IN3(n1106), .QN(n1246));
   NAND4X0 U1186 (.IN1(n1107), .IN2(round[1]), .IN3(round[2]), .IN4(n175), .QN(n1106));
   AO22X1 U1187 (.IN1(round[2]), .IN2(n1108), .IN3(n1109), .IN4(n1107), .Q(n1247));
   AO21X1 U1188 (.IN1(enc_ctrl_reg[0]), .IN2(n177), .IN3(n1110), .Q(n1108));
   AO22X1 U1189 (.IN1(round[1]), .IN2(n1110), .IN3(n1107), .IN4(n177), .Q(n1248));
   AO21X1 U1190 (.IN1(enc_ctrl_reg[0]), .IN2(n178), .IN3(n1111), .Q(n1110));
   AO22X1 U1191 (.IN1(n1111), .IN2(round[0]), .IN3(enc_ctrl_reg[0]), .IN4(n178), .Q(n1249)
          );
   AO21X1 U1192 (.IN1(n1103), .IN2(n1092), .IN3(n1319), .Q(n1250));
   AO21X1 U1194 (.IN1(enc_ctrl_reg[1]), .IN2(n158), .IN3(n1099), .Q(n1251));
   OAI22X1 U1197 (.IN1(n179), .IN2(n1320), .IN3(enc_ctrl_reg[0]), .IN4(n1114), .QN(n1252)
          );
   AOI21X1 U1198 (.IN1(n1320), .IN2(n700), .IN3(n896), .QN(n1114));
   AO22X1 U1199 (.IN1(n1115), .IN2(sword_ctr_reg[0]), .IN3(n1116), .IN4(n1320), .Q(n1253)
          );
   SDFFARX1 \enc_ctrl_reg_reg[0]  (.D(n1250), .SI(n1324), .SE(test_se), .CLK(clk), .RSTB(
          n1267), .Q(enc_ctrl_reg[0]), .QN(n158));
   NAND2X1 U140 (.IN1(n697), .IN2(n895), .QN(n1));
   NAND2X1 U141 (.IN1(n697), .IN2(n698), .QN(n2));
   NAND2X1 U142 (.IN1(n697), .IN2(n1091), .QN(n3));
   NAND2X1 U143 (.IN1(n697), .IN2(n1098), .QN(n4));
   INVX0 U144 (.INP(n895), .ZN(n622));
   INVX0 U145 (.INP(n895), .ZN(n629));
   INVX0 U146 (.INP(n698), .ZN(n483));
   INVX0 U147 (.INP(n698), .ZN(n453));
   INVX0 U148 (.INP(n1091), .ZN(n501));
   INVX0 U149 (.INP(n1091), .ZN(n503));
   INVX0 U150 (.INP(n307), .ZN(n440));
   NBUFFX2 U151 (.INP(n1279), .Z(n1277));
   NBUFFX2 U152 (.INP(n1279), .Z(n1276));
   NBUFFX2 U153 (.INP(n1280), .Z(n1275));
   NBUFFX2 U154 (.INP(n1280), .Z(n1274));
   NBUFFX2 U155 (.INP(n1280), .Z(n1273));
   NBUFFX2 U156 (.INP(n1281), .Z(n1271));
   NBUFFX2 U157 (.INP(n1281), .Z(n1270));
   NBUFFX2 U158 (.INP(n1282), .Z(n1269));
   NBUFFX2 U159 (.INP(n1282), .Z(n1268));
   NBUFFX2 U160 (.INP(n1281), .Z(n1272));
   NBUFFX2 U161 (.INP(n1282), .Z(n1267));
   NBUFFX2 U162 (.INP(n1279), .Z(n1278));
   INVX0 U163 (.INP(n308), .ZN(n572));
   INVX0 U164 (.INP(n310), .ZN(n489));
   NAND2X1 U165 (.IN1(n699), .IN2(n309), .QN(n895));
   INVX0 U166 (.INP(n1), .ZN(n690));
   NAND2X1 U167 (.IN1(n699), .IN2(n307), .QN(n698));
   INVX0 U168 (.INP(n2), .ZN(n770));
   INVX0 U169 (.INP(n1), .ZN(n678));
   INVX0 U170 (.INP(n2), .ZN(n701));
   NAND2X1 U171 (.IN1(n699), .IN2(n310), .QN(n1091));
   INVX0 U172 (.INP(n3), .ZN(n642));
   INVX0 U173 (.INP(n3), .ZN(n672));
   INVX0 U174 (.INP(n4), .ZN(n1265));
   INVX0 U175 (.INP(n4), .ZN(n1266));
   INVX0 U176 (.INP(n1098), .ZN(n579));
   INVX0 U177 (.INP(n1098), .ZN(n592));
   INVX0 U178 (.INP(n1264), .ZN(n1262));
   INVX0 U179 (.INP(n1264), .ZN(n1263));
   INVX0 U180 (.INP(n897), .ZN(n888));
   INVX0 U181 (.INP(n966), .ZN(n876));
   INVX0 U182 (.INP(n1254), .ZN(n1084));
   INVX0 U183 (.INP(n1254), .ZN(n1072));
   NBUFFX2 U184 (.INP(reset_n), .Z(n1280));
   NBUFFX2 U185 (.INP(reset_n), .Z(n1279));
   NBUFFX2 U186 (.INP(reset_n), .Z(n1282));
   NBUFFX2 U187 (.INP(reset_n), .Z(n1281));
   INVX0 U188 (.INP(n307), .ZN(n1315));
   INVX0 U189 (.INP(round_key[59]), .ZN(n1303));
   INVX0 U190 (.INP(round_key[95]), .ZN(n1291));
   INVX0 U191 (.INP(round_key[31]), .ZN(n1307));
   INVX0 U192 (.INP(round_key[27]), .ZN(n1311));
   INVX0 U193 (.INP(round_key[91]), .ZN(n1295));
   INVX0 U194 (.INP(round_key[90]), .ZN(n1296));
   INVX0 U195 (.INP(round_key[58]), .ZN(n1304));
   INVX0 U196 (.INP(round_key[26]), .ZN(n1312));
   INVX0 U197 (.INP(round_key[24]), .ZN(n1314));
   INVX0 U198 (.INP(round_key[25]), .ZN(n1313));
   INVX0 U199 (.INP(round_key[89]), .ZN(n1297));
   INVX0 U200 (.INP(round_key[57]), .ZN(n1305));
   INVX0 U201 (.INP(round_key[56]), .ZN(n1306));
   INVX0 U202 (.INP(round_key[88]), .ZN(n1298));
   INVX0 U203 (.INP(round_key[63]), .ZN(n1299));
   INVX0 U204 (.INP(round_key[93]), .ZN(n1293));
   INVX0 U205 (.INP(round_key[29]), .ZN(n1309));
   INVX0 U206 (.INP(round_key[61]), .ZN(n1301));
   INVX0 U207 (.INP(round_key[28]), .ZN(n1310));
   INVX0 U208 (.INP(round_key[62]), .ZN(n1300));
   INVX0 U209 (.INP(round_key[30]), .ZN(n1308));
   INVX0 U210 (.INP(round_key[92]), .ZN(n1294));
   INVX0 U211 (.INP(round_key[94]), .ZN(n1292));
   INVX0 U212 (.INP(round_key[60]), .ZN(n1302));
   INVX0 U348 (.INP(round_key[123]), .ZN(n1287));
   INVX0 U351 (.INP(round_key[122]), .ZN(n1288));
   INVX0 U356 (.INP(round_key[120]), .ZN(n1290));
   INVX0 U359 (.INP(round_key[121]), .ZN(n1289));
   INVX0 U371 (.INP(round_key[127]), .ZN(n1283));
   INVX0 U374 (.INP(round_key[125]), .ZN(n1285));
   INVX0 U380 (.INP(round_key[124]), .ZN(n1286));
   INVX0 U406 (.INP(round_key[126]), .ZN(n1284));
   NAND2X1 U409 (.IN1(n699), .IN2(n308), .QN(n1098));
   INVX0 U414 (.INP(n1102), .ZN(n1321));
   INVX0 U417 (.INP(n1115), .ZN(n1320));
   XOR3X1 U429 (.IN1(n151), .IN2(n142), .IN3(n771), .Q(n769));
   XNOR2X1 U432 (.IN1(round_key[52]), .IN2(new_block[68]), .Q(n142));
   XOR3X1 U464 (.IN1(n147), .IN2(n143), .IN3(n1067), .Q(n1065));
   XNOR2X1 U468 (.IN1(round_key[4]), .IN2(new_block[76]), .Q(n143));
   XOR3X1 U473 (.IN1(n271), .IN2(n144), .IN3(n454), .Q(n452));
   XNOR2X1 U477 (.IN1(round_key[105]), .IN2(new_block[81]), .Q(n144));
   XOR3X1 U489 (.IN1(n244), .IN2(n145), .IN3(n1073), .Q(n1071));
   XNOR2X1 U492 (.IN1(round_key[3]), .IN2(new_block[75]), .Q(n145));
   XOR3X1 U566 (.IN1(n163), .IN2(n146), .IN3(n877), .Q(n875));
   XNOR2X1 U569 (.IN1(round_key[35]), .IN2(new_block[59]), .Q(n146));
   XOR3X1 U574 (.IN1(n147), .IN2(n148), .IN3(n1017), .Q(n1015));
   XNOR2X1 U577 (.IN1(round_key[12]), .IN2(new_block[36]), .Q(n148));
   XOR3X1 U589 (.IN1(n188), .IN2(n149), .IN3(n673), .Q(n671));
   XNOR2X1 U592 (.IN1(round_key[68]), .IN2(new_block[92]), .Q(n149));
   XOR3X1 U624 (.IN1(n162), .IN2(n150), .IN3(n871), .Q(n869));
   XNOR2X1 U627 (.IN1(round_key[36]), .IN2(new_block[60]), .Q(n150));
   XOR3X1 U632 (.IN1(n151), .IN2(n152), .IN3(n821), .Q(n819));
   XNOR2X1 U635 (.IN1(round_key[44]), .IN2(new_block[68]), .Q(n152));
   XOR3X1 U647 (.IN1(n188), .IN2(n153), .IN3(n623), .Q(n621));
   XNOR2X1 U650 (.IN1(round_key[76]), .IN2(new_block[92]), .Q(n153));
   XOR3X1 U662 (.IN1(n265), .IN2(n154), .IN3(n484), .Q(n482));
   XNOR2X1 U682 (.IN1(round_key[100]), .IN2(new_block[84]), .Q(n154));
   XOR3X1 U686 (.IN1(n193), .IN2(n155), .IN3(n490), .Q(n488));
   XNOR2X1 U691 (.IN1(round_key[99]), .IN2(new_block[83]), .Q(n155));
   XOR3X1 U695 (.IN1(n200), .IN2(n156), .IN3(n967), .Q(n965));
   XNOR2X1 U707 (.IN1(round_key[20]), .IN2(new_block[76]), .Q(n156));
   XOR3X1 U710 (.IN1(n176), .IN2(n205), .IN3(n573), .Q(n571));
   XNOR2X1 U719 (.IN1(round_key[84]), .IN2(new_block[92]), .Q(n205));
   XOR3X1 U792 (.IN1(n165), .IN2(n212), .IN3(n889), .Q(n887));
   XNOR2X1 U795 (.IN1(round_key[33]), .IN2(new_block[57]), .Q(n212));
   XOR3X1 U800 (.IN1(n195), .IN2(n222), .IN3(n502), .Q(n500));
   XNOR2X1 U803 (.IN1(round_key[97]), .IN2(new_block[81]), .Q(n222));
   XOR3X1 U815 (.IN1(n252), .IN2(n242), .IN3(n643), .Q(n641));
   XNOR2X1 U818 (.IN1(round_key[73]), .IN2(new_block[97]), .Q(n242));
   XOR3X1 U830 (.IN1(n250), .IN2(n243), .IN3(n1085), .Q(n1083));
   XNOR2X1 U850 (.IN1(round_key[1]), .IN2(new_block[73]), .Q(n243));
   XOR3X1 U853 (.IN1(n244), .IN2(n245), .IN3(n1024), .Q(n1022));
   XNOR2X1 U858 (.IN1(round_key[11]), .IN2(new_block[35]), .Q(n245));
   XOR3X1 U861 (.IN1(n189), .IN2(n246), .IN3(n679), .Q(n677));
   XNOR2X1 U873 (.IN1(round_key[67]), .IN2(new_block[91]), .Q(n246));
   XOR3X1 U876 (.IN1(n256), .IN2(n247), .IN3(n630), .Q(n628));
   XNOR2X1 U908 (.IN1(round_key[75]), .IN2(new_block[99]), .Q(n247));
   XOR3X1 U912 (.IN1(n203), .IN2(n248), .IN3(n987), .Q(n985));
   XNOR2X1 U917 (.IN1(round_key[17]), .IN2(new_block[73]), .Q(n248));
   XOR3X1 U921 (.IN1(n258), .IN2(n249), .IN3(n828), .Q(n826));
   XNOR2X1 U933 (.IN1(round_key[43]), .IN2(new_block[67]), .Q(n249));
   XOR3X1 U936 (.IN1(n250), .IN2(n251), .IN3(n1037), .Q(n1035));
   XNOR2X1 U945 (.IN1(round_key[9]), .IN2(new_block[33]), .Q(n251));
   XOR3X1 U1018 (.IN1(n252), .IN2(n253), .IN3(n691), .Q(n689));
   XNOR2X1 U1021 (.IN1(round_key[65]), .IN2(new_block[9]), .Q(n253));
   XOR3X1 U1026 (.IN1(n260), .IN2(n254), .IN3(n841), .Q(n839));
   XNOR2X1 U1029 (.IN1(round_key[41]), .IN2(new_block[65]), .Q(n254));
   XOR3X1 U1041 (.IN1(n201), .IN2(n255), .IN3(n974), .Q(n972));
   XNOR2X1 U1044 (.IN1(round_key[19]), .IN2(new_block[75]), .Q(n255));
   XOR3X1 U1076 (.IN1(n256), .IN2(n257), .IN3(n580), .Q(n578));
   XNOR2X1 U1079 (.IN1(round_key[83]), .IN2(new_block[99]), .Q(n257));
   XOR3X1 U1084 (.IN1(n258), .IN2(n259), .IN3(n778), .Q(n776));
   XNOR2X1 U1087 (.IN1(round_key[51]), .IN2(new_block[67]), .Q(n259));
   XOR3X1 U1099 (.IN1(n260), .IN2(n261), .IN3(n791), .Q(n789));
   XNOR2X1 U1102 (.IN1(round_key[49]), .IN2(new_block[65]), .Q(n261));
   XOR3X1 U1134 (.IN1(n262), .IN2(n263), .IN3(n593), .Q(n591));
   XNOR2X1 U1138 (.IN1(round_key[81]), .IN2(new_block[9]), .Q(n263));
   XOR3X1 U1143 (.IN1(n173), .IN2(n264), .IN3(n441), .Q(n439));
   XNOR2X1 U1147 (.IN1(round_key[107]), .IN2(new_block[83]), .Q(n264));
   XOR3X1 U1159 (.IN1(n265), .IN2(n266), .IN3(n384), .Q(n382));
   XNOR2X1 U1162 (.IN1(round_key[116]), .IN2(new_block[4]), .Q(n266));
   XOR3X1 U1171 (.IN1(n172), .IN2(n267), .IN3(n434), .Q(n432));
   XNOR2X1 U1179 (.IN1(round_key[108]), .IN2(new_block[84]), .Q(n267));
   XOR3X1 U1180 (.IN1(round_key[71]), .IN2(n268), .IN3(new_block[94]), .Q(n655));
   XOR3X1 U1193 (.IN1(round_key[47]), .IN2(n269), .IN3(new_block[70]), .Q(n803));
   XOR3X1 U1195 (.IN1(n173), .IN2(n270), .IN3(n391), .Q(n389));
   XNOR2X1 U1196 (.IN1(round_key[115]), .IN2(new_block[43]), .Q(n270));
   XOR3X1 U1200 (.IN1(n271), .IN2(n272), .IN3(n404), .Q(n402));
   XNOR2X1 U1201 (.IN1(round_key[113]), .IN2(new_block[41]), .Q(n272));
   XOR3X1 U1202 (.IN1(round_key[112]), .IN2(n273), .IN3(new_block[120]), .Q(n410));
   NAND3X0 U1203 (.IN1(n180), .IN2(n179), .IN3(n697), .QN(n308));
   OAI22X1 U1204 (.IN1(n177), .IN2(keylen), .IN3(n274), .IN4(n311), .QN(n1112));
   AND2X1 U1205 (.IN1(keylen), .IN2(n177), .Q(n311));
   AO22X1 U1206 (.IN1(enc_ctrl_reg[0]), .IN2(n157), .IN3(n1101), .IN4(n1102), .Q(n1099));
   NOR2X0 U1207 (.IN1(n157), .IN2(enc_ctrl_reg[0]), .QN(n1103));
   NOR2X0 U1208 (.IN1(n157), .IN2(n158), .QN(n1101));
   NOR2X0 U1209 (.IN1(n180), .IN2(sword_ctr_reg[1]), .QN(n700));
   NOR2X0 U1210 (.IN1(n179), .IN2(sword_ctr_reg[0]), .QN(n896));
   NOR2X0 U1211 (.IN1(n179), .IN2(n180), .QN(n1092));
   NAND3X0 U1212 (.IN1(n158), .IN2(n157), .IN3(next), .QN(n1104));
   OA21X1 U1213 (.IN1(round[2]), .IN2(n158), .IN3(n1318), .Q(n1105));
   INVX0 U1214 (.INP(n1108), .ZN(n1318));
   NOR2X0 U1215 (.IN1(round[2]), .IN2(n177), .QN(n1109));
   NOR2X0 U1216 (.IN1(n1103), .IN2(enc_ctrl_reg[0]), .QN(n1115));
   NOR2X0 U1217 (.IN1(sword_ctr_reg[0]), .IN2(enc_ctrl_reg[0]), .QN(n1116));
   NOR2X0 U1218 (.IN1(n178), .IN2(n158), .QN(n1107));
   INVX0 U1219 (.INP(n316), .ZN(n1264));
   INVX0 U1220 (.INP(n1262), .ZN(n1261));
   INVX0 U1221 (.INP(n1263), .ZN(n1256));
   INVX0 U1222 (.INP(n1262), .ZN(n1259));
   INVX0 U1223 (.INP(n1262), .ZN(n1260));
   INVX0 U1224 (.INP(n1263), .ZN(n1258));
   INVX0 U1225 (.INP(n1263), .ZN(n1257));
   INVX0 U1226 (.INP(n316), .ZN(n433));
   INVX0 U1227 (.INP(n1263), .ZN(n1255));
   NAND2X0 U1228 (.IN1(n1321), .IN2(n1101), .QN(n317));
   INVX0 U1229 (.INP(n317), .ZN(n1254));
   INVX0 U1230 (.INP(n317), .ZN(n1113));
   INVX0 U1231 (.INP(n1084), .ZN(n973));
   INVX0 U1232 (.INP(n1072), .ZN(n986));
   INVX0 U1233 (.INP(n1072), .ZN(n1066));
   INVX0 U1234 (.INP(n1084), .ZN(n1016));
   INVX0 U1235 (.INP(n1084), .ZN(n1023));
   INVX0 U1236 (.INP(n1072), .ZN(n1036));
   INVX0 U1237 (.INP(n1084), .ZN(n403));
   INVX0 U1238 (.INP(n318), .ZN(n966));
   INVX0 U1239 (.INP(n318), .ZN(n897));
   INVX0 U1240 (.INP(n876), .ZN(n870));
   INVX0 U1241 (.INP(n888), .ZN(n840));
   INVX0 U1242 (.INP(n876), .ZN(n820));
   INVX0 U1243 (.INP(n876), .ZN(n827));
   INVX0 U1244 (.INP(n888), .ZN(n777));
   INVX0 U1245 (.INP(n888), .ZN(n790));
   INVX0 U1246 (.INP(n888), .ZN(n390));
   INVX0 U1247 (.INP(n310), .ZN(n1316));
   INVX0 U1248 (.INP(n309), .ZN(n383));
   NAND2X0 U1249 (.IN1(n1099), .IN2(n1100), .QN(n316));
   NAND2X0 U1250 (.IN1(round[3]), .IN2(n1112), .QN(n1102));
   NAND2X0 U1251 (.IN1(n1317), .IN2(n1099), .QN(n318));
   INVX0 U1252 (.INP(n1100), .ZN(n1317));
   NOR2X0 U1253 (.IN1(n1099), .IN2(n1317), .QN(n697));
   NAND2X0 U1254 (.IN1(n896), .IN2(n697), .QN(n309));
   NAND2X0 U1255 (.IN1(n1092), .IN2(n697), .QN(n310));
   NAND2X0 U1256 (.IN1(n700), .IN2(n697), .QN(n307));
   NOR2X0 U1257 (.IN1(n1319), .IN2(enc_ctrl_reg[0]), .QN(n1111));
   INVX0 U1258 (.INP(n1104), .ZN(n1319));
endmodule

module aes_inv_sbox (sboxw, new_sboxw);
input [31:0] sboxw;
output [31:0] new_sboxw;
wire n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
       n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199
       , n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
       n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226
       , n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
       n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253
       , n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
       n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280
       , n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
       n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307
       , n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
       n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334
       , n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, 
       n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361
       , n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
       n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388
       , n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
       n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415
       , n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, 
       n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442
       , n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, 
       n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469
       , n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
       n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496
       , n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
       n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523
       , n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, 
       n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550
       , n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, 
       n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577
       , n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
       n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604
       , n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
       n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631
       , n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, 
       n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658
       , n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, 
       n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685
       , n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
       n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712
       , n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
       n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739
       , n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, 
       n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766
       , n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, 
       n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793
       , n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
       n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820
       , n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, 
       n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847
       , n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, 
       n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874
       , n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, 
       n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901
       , n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
       n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928
       , n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
       n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955
       , n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, 
       n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982
       , n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, 
       n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, 
       n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019
       , n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
       n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042
       , n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
       n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065
       , n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, 
       n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088
       , n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
       n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111
       , n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
       n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134
       , n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, 
       n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157
       , n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
       n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180
       , n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, 
       n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203
       , n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
       n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226
       , n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, 
       n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249
       , n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, 
       n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272
       , n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
       n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295
       , n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
       n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318
       , n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
       n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341
       , n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
       n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364
       , n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
       n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387
       , n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
       n1399, n1400, n1401, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
       n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
       , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
       n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64
       , n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, 
       n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
       , n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111
       , n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
       n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138
       , n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
       n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165
       , n166, n167, n168, n169, n170, n171, n1402, n1403, n1404, n1405, n1406, n1407, 
       n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415;
   AO222X1 U678 (.IN1(n172), .IN2(n173), .IN3(n174), .IN4(n175), .IN5(n176), .IN6(n66), .Q(
          new_sboxw[9]));
   AO221X1 U679 (.IN1(n177), .IN2(n178), .IN3(n179), .IN4(n180), .IN5(n181), .Q(n176));
   AO22X1 U680 (.IN1(n182), .IN2(n183), .IN3(n184), .IN4(n185), .Q(n181));
   OA221X1 U681 (.IN1(n188), .IN2(n33), .IN3(n1412), .IN4(n56), .IN5(n189), .Q(n187));
   OA222X1 U682 (.IN1(n60), .IN2(n1411), .IN3(n1409), .IN4(n58), .IN5(n6), .IN6(n43), .Q(
          n186));
   NAND4X0 U683 (.IN1(n190), .IN2(n47), .IN3(n191), .IN4(n192), .QN(n183));
   OA222X1 U684 (.IN1(n193), .IN2(n46), .IN3(n1409), .IN4(n34), .IN5(n194), .IN6(n38), .Q(
          n192));
   NAND4X0 U685 (.IN1(n197), .IN2(n47), .IN3(n198), .IN4(n199), .QN(n180));
   OA222X1 U686 (.IN1(sboxw[11]), .IN2(n1), .IN3(n200), .IN4(n1412), .IN5(n194), .IN6(n35)
          , .Q(n199));
   NAND4X0 U687 (.IN1(n202), .IN2(n196), .IN3(n203), .IN4(n204), .QN(n178));
   OA222X1 U688 (.IN1(n193), .IN2(n43), .IN3(n37), .IN4(n1410), .IN5(n47), .IN6(n1411), .Q(
          n204));
   AO222X1 U689 (.IN1(n205), .IN2(n206), .IN3(n8), .IN4(n207), .IN5(n208), .IN6(n64), .Q(
          n175));
   NAND4X0 U690 (.IN1(n209), .IN2(n210), .IN3(n211), .IN4(n212), .QN(n208));
   OA221X1 U691 (.IN1(n6), .IN2(n213), .IN3(n51), .IN4(n1410), .IN5(n214), .Q(n212));
   NAND4X0 U692 (.IN1(n40), .IN2(n216), .IN3(n217), .IN4(n218), .QN(n207));
   OA22X1 U693 (.IN1(n193), .IN2(n57), .IN3(n219), .IN4(n213), .Q(n218));
   AO221X1 U694 (.IN1(n220), .IN2(n64), .IN3(n221), .IN4(n206), .IN5(n222), .Q(n173));
   OAI21X1 U695 (.IN1(n223), .IN2(n64), .IN3(n224), .QN(n222));
   OA221X1 U696 (.IN1(n219), .IN2(n60), .IN3(n225), .IN4(n46), .IN5(n226), .Q(n223));
   NAND4X0 U697 (.IN1(n45), .IN2(n227), .IN3(n228), .IN4(n229), .QN(n220));
   OA22X1 U698 (.IN1(n1415), .IN2(n43), .IN3(n60), .IN4(n1414), .Q(n229));
   AO21X1 U699 (.IN1(n42), .IN2(n53), .IN3(n1410), .Q(n228));
   AO222X1 U700 (.IN1(n172), .IN2(n230), .IN3(n174), .IN4(n231), .IN5(n232), .IN6(n66), .Q(
          new_sboxw[8]));
   AO222X1 U701 (.IN1(n182), .IN2(n233), .IN3(n184), .IN4(n234), .IN5(sboxw[14]), .IN6(
          n235), .Q(n232));
   AO222X1 U702 (.IN1(n8), .IN2(n236), .IN3(n237), .IN4(n64), .IN5(n238), .IN6(n6), .Q(
          n235));
   AO22X1 U703 (.IN1(n239), .IN2(n1415), .IN3(n240), .IN4(n1411), .Q(n237));
   NAND4X0 U704 (.IN1(n241), .IN2(n43), .IN3(n242), .IN4(n243), .QN(n236));
   OA222X1 U705 (.IN1(n213), .IN2(n1410), .IN3(n219), .IN4(n58), .IN5(n1414), .IN6(n61), .
          Q(n243));
   OR2X1 U706 (.IN1(n244), .IN2(n225), .Q(n242));
   NAND4X0 U707 (.IN1(n245), .IN2(n246), .IN3(n247), .IN4(n248), .QN(n234));
   OR2X1 U708 (.IN1(n1414), .IN2(n249), .Q(n247));
   NAND3X0 U709 (.IN1(n252), .IN2(n244), .IN3(n253), .QN(n233));
   OA221X1 U710 (.IN1(n6), .IN2(n57), .IN3(n254), .IN4(n1), .IN5(n209), .Q(n253));
   OA22X1 U711 (.IN1(n1412), .IN2(n53), .IN3(n225), .IN4(n60), .Q(n252));
   NAND3X0 U712 (.IN1(n255), .IN2(n256), .IN3(n257), .QN(n231));
   OA222X1 U713 (.IN1(n63), .IN2(n46), .IN3(n8), .IN4(n258), .IN5(n259), .IN6(n64), .Q(
          n257));
   OA221X1 U714 (.IN1(n219), .IN2(n61), .IN3(n1409), .IN4(n58), .IN5(n260), .Q(n259));
   OA221X1 U715 (.IN1(n194), .IN2(n53), .IN3(n225), .IN4(n58), .IN5(n263), .Q(n258));
   AND2X1 U716 (.IN1(n47), .IN2(n264), .Q(n263));
   AO221X1 U717 (.IN1(n265), .IN2(n64), .IN3(n8), .IN4(n266), .IN5(n267), .Q(n230));
   AO22X1 U718 (.IN1(n206), .IN2(n268), .IN3(n269), .IN4(n1414), .Q(n267));
   NAND4X0 U719 (.IN1(n270), .IN2(n38), .IN3(n271), .IN4(n272), .QN(n266));
   OA22X1 U720 (.IN1(n225), .IN2(n57), .IN3(n1415), .IN4(n53), .Q(n272));
   AO221X1 U721 (.IN1(n225), .IN2(n273), .IN3(n261), .IN4(n1413), .IN5(n274), .Q(n265));
   AO21X1 U722 (.IN1(n53), .IN2(n35), .IN3(n219), .Q(n275));
   AO22X1 U723 (.IN1(n276), .IN2(n1408), .IN3(sboxw[7]), .IN4(n277), .Q(new_sboxw[7]));
   AO22X1 U724 (.IN1(n278), .IN2(n1407), .IN3(sboxw[6]), .IN4(n279), .Q(n277));
   AO222X1 U725 (.IN1(n280), .IN2(n281), .IN3(n13), .IN4(n282), .IN5(n283), .IN6(n14), .Q(
          n279));
   NAND4X0 U726 (.IN1(n284), .IN2(n285), .IN3(n286), .IN4(n287), .QN(n283));
   AO221X1 U727 (.IN1(n155), .IN2(n27), .IN3(n291), .IN4(n25), .IN5(n292), .Q(n282));
   NAND4X0 U728 (.IN1(n293), .IN2(n294), .IN3(n295), .IN4(n296), .QN(n278));
   OA221X1 U729 (.IN1(n297), .IN2(n1404), .IN3(n107), .IN4(n154), .IN5(n298), .Q(n296));
   NAND4X0 U730 (.IN1(n28), .IN2(n152), .IN3(n300), .IN4(n301), .QN(n299));
   OA22X1 U731 (.IN1(n5), .IN2(n165), .IN3(n302), .IN4(n154), .Q(n301));
   AO221X1 U732 (.IN1(n305), .IN2(n4), .IN3(n306), .IN4(n27), .IN5(n307), .Q(n304));
   AO222X1 U733 (.IN1(n308), .IN2(n309), .IN3(n310), .IN4(n311), .IN5(sboxw[6]), .IN6(n312)
          , .Q(n276));
   AO221X1 U734 (.IN1(n313), .IN2(n14), .IN3(n303), .IN4(n281), .IN5(n314), .Q(n312));
   AO21X1 U735 (.IN1(n13), .IN2(n315), .IN3(n316), .Q(n314));
   AO221X1 U736 (.IN1(n317), .IN2(n22), .IN3(n318), .IN4(n319), .IN5(n320), .Q(n315));
   NAND4X0 U737 (.IN1(n321), .IN2(n160), .IN3(n322), .IN4(n323), .QN(n313));
   OA22X1 U738 (.IN1(n4), .IN2(n151), .IN3(n288), .IN4(n164), .Q(n323));
   NAND4X0 U739 (.IN1(n324), .IN2(n325), .IN3(n326), .IN4(n327), .QN(n311));
   OA22X1 U740 (.IN1(n5), .IN2(n162), .IN3(n288), .IN4(n159), .Q(n327));
   AO221X1 U741 (.IN1(n328), .IN2(n329), .IN3(n330), .IN4(n302), .IN5(n331), .Q(n309));
   AO221X1 U742 (.IN1(n332), .IN2(n25), .IN3(n333), .IN4(n334), .IN5(n335), .Q(n331));
   AO222X1 U743 (.IN1(n336), .IN2(n337), .IN3(n338), .IN4(n339), .IN5(sboxw[7]), .IN6(n340)
          , .Q(new_sboxw[6]));
   AO222X1 U744 (.IN1(n310), .IN2(n341), .IN3(sboxw[6]), .IN4(n342), .IN5(n308), .IN6(n343)
          , .Q(n340));
   NAND4X0 U745 (.IN1(n344), .IN2(n345), .IN3(n346), .IN4(n347), .QN(n343));
   OA221X1 U746 (.IN1(n1404), .IN2(n22), .IN3(n165), .IN4(n29), .IN5(n348), .Q(n347));
   OA22X1 U747 (.IN1(n30), .IN2(n151), .IN3(n328), .IN4(n156), .Q(n346));
   AO22X1 U748 (.IN1(n13), .IN2(n349), .IN3(n350), .IN4(n14), .Q(n342));
   NAND4X0 U749 (.IN1(n351), .IN2(n352), .IN3(n353), .IN4(n354), .QN(n350));
   OA222X1 U750 (.IN1(n355), .IN2(n1405), .IN3(n27), .IN4(n157), .IN5(n152), .IN6(n22), .Q(
          n354));
   AND2X1 U751 (.IN1(n356), .IN2(n357), .Q(n353));
   NAND4X0 U752 (.IN1(n358), .IN2(n359), .IN3(n360), .IN4(n361), .QN(n349));
   AND4X1 U753 (.IN1(n345), .IN2(n362), .IN3(n363), .IN4(n357), .Q(n361));
   OA22X1 U754 (.IN1(n25), .IN2(n1402), .IN3(n5), .IN4(n152), .Q(n360));
   NAND4X0 U755 (.IN1(n357), .IN2(n325), .IN3(n365), .IN4(n366), .QN(n341));
   OA22X1 U756 (.IN1(n334), .IN2(n160), .IN3(n319), .IN4(n171), .Q(n366));
   AO22X1 U757 (.IN1(n13), .IN2(n367), .IN3(n368), .IN4(n14), .Q(n339));
   NAND4X0 U758 (.IN1(n294), .IN2(n157), .IN3(n369), .IN4(n370), .QN(n368));
   OA222X1 U759 (.IN1(n319), .IN2(n159), .IN3(n5), .IN4(n165), .IN5(n328), .IN6(n164), .Q(
          n370));
   OA22X1 U760 (.IN1(n160), .IN2(n29), .IN3(n106), .IN4(n171), .Q(n369));
   NAND4X0 U761 (.IN1(n345), .IN2(n158), .IN3(n21), .IN4(n371), .QN(n367));
   OA222X1 U762 (.IN1(n4), .IN2(n159), .IN3(n5), .IN4(n167), .IN5(n25), .IN6(n151), .Q(
          n371));
   NAND3X0 U763 (.IN1(n351), .IN2(n372), .IN3(n373), .QN(n337));
   OA22X1 U764 (.IN1(n374), .IN2(n14), .IN3(n13), .IN4(n375), .Q(n373));
   OA221X1 U765 (.IN1(n1404), .IN2(n25), .IN3(n5), .IN4(n158), .IN5(n376), .Q(n375));
   OA22X1 U766 (.IN1(n302), .IN2(n1405), .IN3(sboxw[2]), .IN4(n328), .Q(n376));
   OA221X1 U767 (.IN1(n355), .IN2(n1402), .IN3(n377), .IN4(n30), .IN5(n357), .Q(n374));
   AO222X1 U768 (.IN1(n336), .IN2(n378), .IN3(n338), .IN4(n379), .IN5(sboxw[7]), .IN6(n380)
          , .Q(new_sboxw[5]));
   AO221X1 U769 (.IN1(n310), .IN2(n381), .IN3(n308), .IN4(n382), .IN5(n383), .Q(n380));
   AO22X1 U770 (.IN1(n384), .IN2(n385), .IN3(n386), .IN4(n387), .Q(n383));
   NAND4X0 U771 (.IN1(n388), .IN2(n285), .IN3(n389), .IN4(n390), .QN(n387));
   OA222X1 U772 (.IN1(n334), .IN2(n153), .IN3(n25), .IN4(n154), .IN5(n106), .IN6(n164), .Q(
          n390));
   OA22X1 U773 (.IN1(n391), .IN2(n22), .IN3(n4), .IN4(n158), .Q(n389));
   NAND3X0 U774 (.IN1(n348), .IN2(n392), .IN3(n393), .QN(n385));
   OA221X1 U775 (.IN1(n334), .IN2(n1404), .IN3(n5), .IN4(n394), .IN5(n395), .Q(n393));
   NAND3X0 U776 (.IN1(n396), .IN2(n397), .IN3(n398), .QN(n382));
   OA221X1 U777 (.IN1(n319), .IN2(n166), .IN3(n399), .IN4(n27), .IN5(n400), .Q(n398));
   OA22X1 U778 (.IN1(n30), .IN2(n164), .IN3(n401), .IN4(n25), .Q(n396));
   NAND4X0 U779 (.IN1(n20), .IN2(n362), .IN3(n402), .IN4(n403), .QN(n381));
   OA222X1 U780 (.IN1(n334), .IN2(n152), .IN3(n162), .IN4(n25), .IN5(n106), .IN6(n154), .Q(
          n403));
   AO22X1 U781 (.IN1(n13), .IN2(n406), .IN3(n407), .IN4(n14), .Q(n379));
   NAND4X0 U782 (.IN1(n408), .IN2(n409), .IN3(n410), .IN4(n411), .QN(n407));
   AND4X1 U783 (.IN1(n162), .IN2(n325), .IN3(n28), .IN4(n412), .Q(n411));
   OA22X1 U784 (.IN1(n288), .IN2(n151), .IN3(n27), .IN4(n156), .Q(n410));
   NAND4X0 U785 (.IN1(n405), .IN2(n31), .IN3(n414), .IN4(n415), .QN(n406));
   OA222X1 U786 (.IN1(n4), .IN2(n153), .IN3(n328), .IN4(n151), .IN5(n25), .IN6(n158), .Q(
          n415));
   AND2X1 U787 (.IN1(n362), .IN2(n285), .Q(n414));
   AO221X1 U788 (.IN1(n303), .IN2(n281), .IN3(n416), .IN4(n24), .IN5(n417), .Q(n378));
   AO221X1 U789 (.IN1(n13), .IN2(n418), .IN3(n419), .IN4(n14), .IN5(n23), .Q(n417));
   NAND3X0 U790 (.IN1(n334), .IN2(n13), .IN3(n420), .QN(n372));
   NAND4X0 U791 (.IN1(n359), .IN2(n164), .IN3(n421), .IN4(n422), .QN(n419));
   AO222X1 U792 (.IN1(n336), .IN2(n426), .IN3(n338), .IN4(n427), .IN5(sboxw[7]), .IN6(n428)
          , .Q(new_sboxw[4]));
   AO221X1 U793 (.IN1(n386), .IN2(n429), .IN3(n384), .IN4(n430), .IN5(n431), .Q(n428));
   AO22X1 U794 (.IN1(n308), .IN2(n432), .IN3(n310), .IN4(n433), .Q(n431));
   NAND4X0 U795 (.IN1(n294), .IN2(n363), .IN3(n412), .IN4(n434), .QN(n433));
   AOI222X1 U796 (.IN1(n319), .IN2(n291), .IN3(n30), .IN4(n435), .IN5(n305), .IN6(n425), .
          QN(n434));
   NAND4X0 U797 (.IN1(n436), .IN2(n356), .IN3(n437), .IN4(n438), .QN(n432));
   OA222X1 U798 (.IN1(n5), .IN2(n152), .IN3(n302), .IN4(n158), .IN5(n334), .IN6(n157), .Q(
          n438));
   NAND4X0 U799 (.IN1(n405), .IN2(n440), .IN3(n441), .IN4(n442), .QN(n430));
   OA221X1 U800 (.IN1(n106), .IN2(n162), .IN3(n165), .IN4(n26), .IN5(n423), .Q(n442));
   AO21X1 U801 (.IN1(n153), .IN2(n164), .IN3(n29), .Q(n441));
   OA221X1 U802 (.IN1(n288), .IN2(n165), .IN3(n302), .IN4(n167), .IN5(n395), .Q(n444));
   OA222X1 U803 (.IN1(n401), .IN2(n106), .IN3(n4), .IN4(n157), .IN5(n5), .IN6(n154), .Q(
          n443));
   AO222X1 U804 (.IN1(n445), .IN2(n14), .IN3(n13), .IN4(n446), .IN5(n281), .IN6(n307), .Q(
          n427));
   NAND4X0 U805 (.IN1(n28), .IN2(n164), .IN3(n324), .IN4(n447), .QN(n446));
   OA22X1 U806 (.IN1(n425), .IN2(n1402), .IN3(n162), .IN4(n22), .Q(n447));
   NAND4X0 U807 (.IN1(n448), .IN2(n449), .IN3(n450), .IN4(n451), .QN(n445));
   OA222X1 U808 (.IN1(n4), .IN2(n1405), .IN3(n25), .IN4(n157), .IN5(n164), .IN6(n26), .Q(
          n451));
   AO222X1 U809 (.IN1(n281), .IN2(n435), .IN3(n13), .IN4(n452), .IN5(n453), .IN6(n14), .Q(
          n426));
   NAND4X0 U810 (.IN1(n28), .IN2(n436), .IN3(n454), .IN4(n455), .QN(n453));
   OA221X1 U811 (.IN1(n106), .IN2(n162), .IN3(n328), .IN4(n456), .IN5(n457), .Q(n455));
   AND2X1 U812 (.IN1(n345), .IN2(n325), .Q(n454));
   NAND4X0 U813 (.IN1(n458), .IN2(n325), .IN3(n439), .IN4(n459), .QN(n452));
   OA22X1 U814 (.IN1(n425), .IN2(n171), .IN3(n25), .IN4(n154), .Q(n459));
   OA22X1 U815 (.IN1(n29), .IN2(sboxw[2]), .IN3(n25), .IN4(n163), .Q(n425));
   AO22X1 U816 (.IN1(sboxw[7]), .IN2(n460), .IN3(n461), .IN4(n1408), .Q(new_sboxw[3]));
   AO222X1 U817 (.IN1(n384), .IN2(n462), .IN3(n386), .IN4(n463), .IN5(n464), .IN6(n1407), .
          Q(n461));
   AO222X1 U818 (.IN1(n281), .IN2(n161), .IN3(n13), .IN4(n465), .IN5(n466), .IN6(n14), .Q(
          n464));
   NAND4X0 U819 (.IN1(n467), .IN2(n439), .IN3(n468), .IN4(n469), .QN(n466));
   AND3X1 U820 (.IN1(n344), .IN2(n395), .IN3(n448), .Q(n469));
   NAND4X0 U821 (.IN1(n471), .IN2(n321), .IN3(n18), .IN4(n395), .QN(n465));
   OR2X1 U822 (.IN1(n25), .IN2(n289), .Q(n471));
   NAND4X0 U823 (.IN1(n440), .IN2(n154), .IN3(n351), .IN4(n473), .QN(n463));
   OA222X1 U824 (.IN1(n4), .IN2(n1405), .IN3(n288), .IN4(n474), .IN5(n397), .IN6(n30), .Q(
          n473));
   NAND4X0 U825 (.IN1(n477), .IN2(n449), .IN3(n478), .IN4(n479), .QN(n462));
   OA221X1 U826 (.IN1(n152), .IN2(n29), .IN3(n30), .IN4(n158), .IN5(n468), .Q(n479));
   AND2X1 U827 (.IN1(n356), .IN2(n31), .Q(n478));
   AO222X1 U828 (.IN1(n308), .IN2(n481), .IN3(n310), .IN4(n482), .IN5(sboxw[6]), .IN6(n483)
          , .Q(n460));
   AO222X1 U829 (.IN1(n281), .IN2(n291), .IN3(n13), .IN4(n484), .IN5(n485), .IN6(n14), .Q(
          n483));
   NAND4X0 U830 (.IN1(n436), .IN2(n344), .IN3(n486), .IN4(n487), .QN(n485));
   OA222X1 U831 (.IN1(n30), .IN2(n162), .IN3(n404), .IN4(n106), .IN5(n22), .IN6(n1402), .Q(
          n487));
   AO21X1 U832 (.IN1(n153), .IN2(n154), .IN3(n328), .Q(n486));
   NAND4X0 U833 (.IN1(n477), .IN2(n457), .IN3(n488), .IN4(n489), .QN(n484));
   OA221X1 U834 (.IN1(n401), .IN2(n25), .IN3(n159), .IN4(n29), .IN5(n490), .Q(n489));
   NAND4X0 U835 (.IN1(n388), .IN2(n345), .IN3(n491), .IN4(n492), .QN(n482));
   OA222X1 U836 (.IN1(n334), .IN2(n159), .IN3(n493), .IN4(n29), .IN5(n302), .IN6(n156), .Q(
          n492));
   NAND4X0 U837 (.IN1(n18), .IN2(n440), .IN3(n424), .IN4(n494), .QN(n481));
   OA22X1 U838 (.IN1(n328), .IN2(n391), .IN3(n30), .IN4(n164), .Q(n494));
   AO22X1 U839 (.IN1(n496), .IN2(n170), .IN3(sboxw[31]), .IN4(n497), .Q(new_sboxw[31]));
   AO22X1 U840 (.IN1(n498), .IN2(n169), .IN3(sboxw[30]), .IN4(n499), .Q(n497));
   AO222X1 U841 (.IN1(n500), .IN2(n501), .IN3(n3), .IN4(n502), .IN5(n503), .IN6(n17), .Q(
          n499));
   NAND4X0 U842 (.IN1(n504), .IN2(n505), .IN3(n506), .IN4(n507), .QN(n503));
   AO221X1 U843 (.IN1(n131), .IN2(n120), .IN3(n511), .IN4(n118), .IN5(n512), .Q(n502));
   NAND4X0 U844 (.IN1(n513), .IN2(n514), .IN3(n515), .IN4(n516), .QN(n498));
   OA221X1 U845 (.IN1(n517), .IN2(n148), .IN3(n126), .IN4(n130), .IN5(n518), .Q(n516));
   NAND4X0 U846 (.IN1(n121), .IN2(n128), .IN3(n520), .IN4(n521), .QN(n519));
   OA22X1 U847 (.IN1(n12), .IN2(n141), .IN3(n522), .IN4(n130), .Q(n521));
   AO221X1 U848 (.IN1(n525), .IN2(n11), .IN3(n526), .IN4(n120), .IN5(n527), .Q(n524));
   AO222X1 U849 (.IN1(n528), .IN2(n529), .IN3(n530), .IN4(n531), .IN5(sboxw[30]), .IN6(
          n532), .Q(n496));
   AO221X1 U850 (.IN1(n533), .IN2(n17), .IN3(n523), .IN4(n501), .IN5(n534), .Q(n532));
   AO21X1 U851 (.IN1(n3), .IN2(n535), .IN3(n536), .Q(n534));
   AO221X1 U852 (.IN1(n537), .IN2(n115), .IN3(n538), .IN4(n539), .IN5(n540), .Q(n535));
   NAND4X0 U853 (.IN1(n541), .IN2(n136), .IN3(n542), .IN4(n543), .QN(n533));
   OA22X1 U854 (.IN1(n11), .IN2(n127), .IN3(n508), .IN4(n140), .Q(n543));
   NAND4X0 U855 (.IN1(n544), .IN2(n545), .IN3(n546), .IN4(n547), .QN(n531));
   OA22X1 U856 (.IN1(n12), .IN2(n138), .IN3(n508), .IN4(n135), .Q(n547));
   AO221X1 U857 (.IN1(n548), .IN2(n549), .IN3(n550), .IN4(n522), .IN5(n551), .Q(n529));
   AO221X1 U858 (.IN1(n552), .IN2(n118), .IN3(n553), .IN4(n554), .IN5(n555), .Q(n551));
   AO222X1 U859 (.IN1(n556), .IN2(n557), .IN3(n558), .IN4(n559), .IN5(sboxw[31]), .IN6(
          n560), .Q(new_sboxw[30]));
   AO222X1 U860 (.IN1(n530), .IN2(n561), .IN3(sboxw[30]), .IN4(n562), .IN5(n528), .IN6(
          n563), .Q(n560));
   NAND4X0 U861 (.IN1(n564), .IN2(n565), .IN3(n566), .IN4(n567), .QN(n563));
   OA221X1 U862 (.IN1(n148), .IN2(n115), .IN3(n141), .IN4(n122), .IN5(n568), .Q(n567));
   OA22X1 U863 (.IN1(n123), .IN2(n127), .IN3(n548), .IN4(n132), .Q(n566));
   AO22X1 U864 (.IN1(sboxw[29]), .IN2(n569), .IN3(n570), .IN4(n17), .Q(n562));
   NAND4X0 U865 (.IN1(n571), .IN2(n572), .IN3(n573), .IN4(n574), .QN(n570));
   OA222X1 U866 (.IN1(n575), .IN2(n149), .IN3(n120), .IN4(n133), .IN5(n128), .IN6(n115), .
          Q(n574));
   AND2X1 U867 (.IN1(n576), .IN2(n577), .Q(n573));
   NAND4X0 U868 (.IN1(n578), .IN2(n579), .IN3(n580), .IN4(n581), .QN(n569));
   AND4X1 U869 (.IN1(n565), .IN2(n582), .IN3(n583), .IN4(n577), .Q(n581));
   OA22X1 U870 (.IN1(n118), .IN2(n146), .IN3(n12), .IN4(n128), .Q(n580));
   NAND4X0 U871 (.IN1(n577), .IN2(n545), .IN3(n585), .IN4(n586), .QN(n561));
   OA22X1 U872 (.IN1(n554), .IN2(n136), .IN3(n539), .IN4(n145), .Q(n586));
   AO22X1 U873 (.IN1(sboxw[29]), .IN2(n587), .IN3(n588), .IN4(n17), .Q(n559));
   NAND4X0 U874 (.IN1(n514), .IN2(n133), .IN3(n589), .IN4(n590), .QN(n588));
   OA222X1 U875 (.IN1(n539), .IN2(n135), .IN3(n12), .IN4(n141), .IN5(n548), .IN6(n140), .Q(
          n590));
   OA22X1 U876 (.IN1(n136), .IN2(n122), .IN3(n125), .IN4(n145), .Q(n589));
   NAND4X0 U877 (.IN1(n565), .IN2(n134), .IN3(n114), .IN4(n591), .QN(n587));
   OA222X1 U878 (.IN1(n11), .IN2(n135), .IN3(n12), .IN4(n143), .IN5(n118), .IN6(n127), .Q(
          n591));
   NAND3X0 U879 (.IN1(n571), .IN2(n592), .IN3(n593), .QN(n557));
   OA22X1 U880 (.IN1(n594), .IN2(n17), .IN3(n3), .IN4(n595), .Q(n593));
   OA221X1 U881 (.IN1(n148), .IN2(n118), .IN3(n12), .IN4(n134), .IN5(n596), .Q(n595));
   OA22X1 U882 (.IN1(n522), .IN2(n149), .IN3(sboxw[26]), .IN4(n548), .Q(n596));
   OA221X1 U883 (.IN1(n575), .IN2(n146), .IN3(n597), .IN4(n123), .IN5(n577), .Q(n594));
   AO222X1 U884 (.IN1(n598), .IN2(n599), .IN3(n600), .IN4(n601), .IN5(n602), .IN6(n1408), .
          Q(new_sboxw[2]));
   AO222X1 U885 (.IN1(n308), .IN2(n603), .IN3(n310), .IN4(n604), .IN5(sboxw[6]), .IN6(n605)
          , .Q(n602));
   NAND4X0 U886 (.IN1(n321), .IN2(n356), .IN3(n606), .IN4(n607), .QN(n605));
   OA22X1 U887 (.IN1(n13), .IN2(n608), .IN3(n162), .IN4(n107), .Q(n607));
   AO222X1 U888 (.IN1(n288), .IN2(n291), .IN3(n476), .IN4(n106), .IN5(sboxw[3]), .IN6(n22)
          , .Q(n610));
   AO221X1 U889 (.IN1(n329), .IN2(n319), .IN3(n413), .IN4(n5), .IN5(n305), .Q(n609));
   NAND3X0 U890 (.IN1(n31), .IN2(n363), .IN3(n352), .QN(n611));
   NAND4X0 U891 (.IN1(n457), .IN2(n612), .IN3(n613), .IN4(n614), .QN(n604));
   OAI21X1 U892 (.IN1(n152), .IN2(n334), .IN3(n409), .QN(n292));
   OR2X1 U893 (.IN1(n26), .IN2(n391), .Q(n613));
   NAND4X0 U894 (.IN1(n448), .IN2(n458), .IN3(n616), .IN4(n617), .QN(n603));
   OA221X1 U895 (.IN1(n164), .IN2(n22), .IN3(n319), .IN4(n154), .IN5(n298), .Q(n617));
   OA22X1 U896 (.IN1(n158), .IN2(n29), .IN3(n5), .IN4(n157), .Q(n616));
   AO22X1 U897 (.IN1(n13), .IN2(n619), .IN3(n620), .IN4(n14), .Q(n601));
   AO221X1 U898 (.IN1(n618), .IN2(n25), .IN3(n335), .IN4(n26), .IN5(n621), .Q(n620));
   AO221X1 U899 (.IN1(n622), .IN2(n22), .IN3(n302), .IN4(n305), .IN5(n476), .Q(n621));
   NAND4X0 U900 (.IN1(n412), .IN2(n284), .IN3(n623), .IN4(n624), .QN(n619));
   OA222X1 U901 (.IN1(n27), .IN2(n157), .IN3(n493), .IN4(n30), .IN5(n158), .IN6(n29), .Q(
          n624));
   AND2X1 U902 (.IN1(n20), .IN2(n321), .Q(n623));
   AO22X1 U903 (.IN1(n13), .IN2(n626), .IN3(n627), .IN4(n14), .Q(n599));
   NAND4X0 U904 (.IN1(n324), .IN2(n477), .IN3(n628), .IN4(n629), .QN(n627));
   OA222X1 U905 (.IN1(n5), .IN2(n164), .IN3(n328), .IN4(n158), .IN5(n165), .IN6(n29), .Q(
          n629));
   AND2X1 U906 (.IN1(n345), .IN2(n458), .Q(n628));
   NAND4X0 U907 (.IN1(n388), .IN2(n284), .IN3(n630), .IN4(n631), .QN(n626));
   OA222X1 U908 (.IN1(n153), .IN2(n29), .IN3(n328), .IN4(n157), .IN5(n319), .IN6(n154), .Q(
          n631));
   AO222X1 U909 (.IN1(n556), .IN2(n632), .IN3(n558), .IN4(n633), .IN5(sboxw[31]), .IN6(
          n634), .Q(new_sboxw[29]));
   AO221X1 U910 (.IN1(n530), .IN2(n635), .IN3(n528), .IN4(n636), .IN5(n637), .Q(n634));
   AO22X1 U911 (.IN1(n638), .IN2(n639), .IN3(n640), .IN4(n641), .Q(n637));
   NAND4X0 U912 (.IN1(n642), .IN2(n505), .IN3(n643), .IN4(n644), .QN(n641));
   OA222X1 U913 (.IN1(n554), .IN2(n129), .IN3(n118), .IN4(n130), .IN5(n125), .IN6(n140), .
          Q(n644));
   OA22X1 U914 (.IN1(n645), .IN2(n115), .IN3(n11), .IN4(n134), .Q(n643));
   NAND3X0 U915 (.IN1(n568), .IN2(n646), .IN3(n647), .QN(n639));
   OA221X1 U916 (.IN1(n554), .IN2(n148), .IN3(n12), .IN4(n648), .IN5(n649), .Q(n647));
   NAND3X0 U917 (.IN1(n650), .IN2(n651), .IN3(n652), .QN(n636));
   OA221X1 U918 (.IN1(n539), .IN2(n142), .IN3(n653), .IN4(n120), .IN5(n654), .Q(n652));
   OA22X1 U919 (.IN1(n123), .IN2(n140), .IN3(n655), .IN4(n118), .Q(n650));
   NAND4X0 U920 (.IN1(n113), .IN2(n582), .IN3(n656), .IN4(n657), .QN(n635));
   OA222X1 U921 (.IN1(n554), .IN2(n128), .IN3(n138), .IN4(n118), .IN5(n125), .IN6(n130), .
          Q(n657));
   AO22X1 U922 (.IN1(sboxw[29]), .IN2(n660), .IN3(n661), .IN4(n17), .Q(n633));
   NAND4X0 U923 (.IN1(n662), .IN2(n663), .IN3(n664), .IN4(n665), .QN(n661));
   AND4X1 U924 (.IN1(n138), .IN2(n545), .IN3(n121), .IN4(n666), .Q(n665));
   OA22X1 U925 (.IN1(n508), .IN2(n127), .IN3(n120), .IN4(n132), .Q(n664));
   NAND4X0 U926 (.IN1(n659), .IN2(n124), .IN3(n668), .IN4(n669), .QN(n660));
   OA222X1 U927 (.IN1(n11), .IN2(n129), .IN3(n548), .IN4(n127), .IN5(n118), .IN6(n134), .Q(
          n669));
   AND2X1 U928 (.IN1(n582), .IN2(n505), .Q(n668));
   AO221X1 U929 (.IN1(n523), .IN2(n501), .IN3(n670), .IN4(n117), .IN5(n671), .Q(n632));
   NAND4X0 U932 (.IN1(n579), .IN2(n140), .IN3(n675), .IN4(n676), .QN(n673));
   AO222X1 U933 (.IN1(n556), .IN2(n680), .IN3(n558), .IN4(n681), .IN5(sboxw[31]), .IN6(
          n682), .Q(new_sboxw[28]));
   AO221X1 U934 (.IN1(n640), .IN2(n683), .IN3(n638), .IN4(n684), .IN5(n685), .Q(n682));
   AO22X1 U935 (.IN1(n528), .IN2(n686), .IN3(n530), .IN4(n687), .Q(n685));
   NAND4X0 U936 (.IN1(n514), .IN2(n583), .IN3(n666), .IN4(n688), .QN(n687));
   AOI222X1 U937 (.IN1(n539), .IN2(n511), .IN3(n123), .IN4(n689), .IN5(n525), .IN6(n679), .
          QN(n688));
   NAND4X0 U938 (.IN1(n690), .IN2(n576), .IN3(n691), .IN4(n692), .QN(n686));
   OA222X1 U939 (.IN1(n12), .IN2(n128), .IN3(n522), .IN4(n134), .IN5(n554), .IN6(n133), .Q(
          n692));
   NAND4X0 U940 (.IN1(n659), .IN2(n694), .IN3(n695), .IN4(n696), .QN(n684));
   OA221X1 U941 (.IN1(n125), .IN2(n138), .IN3(n141), .IN4(n119), .IN5(n677), .Q(n696));
   AO21X1 U942 (.IN1(n129), .IN2(n140), .IN3(n2), .Q(n695));
   OA221X1 U943 (.IN1(n508), .IN2(n141), .IN3(n522), .IN4(n143), .IN5(n649), .Q(n698));
   OA222X1 U944 (.IN1(n655), .IN2(n125), .IN3(n11), .IN4(n133), .IN5(n12), .IN6(n130), .Q(
          n697));
   AO222X1 U945 (.IN1(n699), .IN2(n17), .IN3(n3), .IN4(n700), .IN5(n501), .IN6(n527), .Q(
          n681));
   NAND4X0 U946 (.IN1(n121), .IN2(n140), .IN3(n544), .IN4(n701), .QN(n700));
   OA22X1 U947 (.IN1(n679), .IN2(n146), .IN3(n138), .IN4(n115), .Q(n701));
   NAND4X0 U948 (.IN1(n702), .IN2(n703), .IN3(n704), .IN4(n705), .QN(n699));
   OA222X1 U949 (.IN1(n11), .IN2(n149), .IN3(n118), .IN4(n133), .IN5(n140), .IN6(n119), .Q(
          n705));
   AO222X1 U950 (.IN1(n501), .IN2(n689), .IN3(n3), .IN4(n706), .IN5(n707), .IN6(n17), .Q(
          n680));
   NAND4X0 U951 (.IN1(n121), .IN2(n690), .IN3(n708), .IN4(n709), .QN(n707));
   OA221X1 U952 (.IN1(n125), .IN2(n138), .IN3(n548), .IN4(n710), .IN5(n711), .Q(n709));
   AND2X1 U953 (.IN1(n565), .IN2(n545), .Q(n708));
   NAND4X0 U954 (.IN1(n712), .IN2(n545), .IN3(n693), .IN4(n713), .QN(n706));
   OA22X1 U955 (.IN1(n679), .IN2(n145), .IN3(n118), .IN4(n130), .Q(n713));
   OA22X1 U956 (.IN1(n2), .IN2(sboxw[26]), .IN3(n118), .IN4(n139), .Q(n679));
   AO22X1 U957 (.IN1(sboxw[31]), .IN2(n714), .IN3(n715), .IN4(n170), .Q(new_sboxw[27]));
   AO222X1 U958 (.IN1(n638), .IN2(n716), .IN3(n640), .IN4(n717), .IN5(n718), .IN6(n169), .
          Q(n715));
   AO222X1 U959 (.IN1(n501), .IN2(n137), .IN3(n3), .IN4(n719), .IN5(n720), .IN6(n17), .Q(
          n718));
   NAND4X0 U960 (.IN1(n721), .IN2(n693), .IN3(n722), .IN4(n723), .QN(n720));
   AND3X1 U961 (.IN1(n564), .IN2(n649), .IN3(n702), .Q(n723));
   NAND4X0 U962 (.IN1(n725), .IN2(n541), .IN3(n111), .IN4(n649), .QN(n719));
   OR2X1 U963 (.IN1(n118), .IN2(n509), .Q(n725));
   NAND4X0 U964 (.IN1(n694), .IN2(n130), .IN3(n571), .IN4(n727), .QN(n717));
   OA222X1 U965 (.IN1(n11), .IN2(n149), .IN3(n508), .IN4(n728), .IN5(n651), .IN6(n123), .Q(
          n727));
   NAND4X0 U966 (.IN1(n731), .IN2(n703), .IN3(n732), .IN4(n733), .QN(n716));
   OA221X1 U967 (.IN1(n128), .IN2(n122), .IN3(n123), .IN4(n134), .IN5(n722), .Q(n733));
   AND2X1 U968 (.IN1(n576), .IN2(n124), .Q(n732));
   AO222X1 U969 (.IN1(n528), .IN2(n735), .IN3(n530), .IN4(n736), .IN5(sboxw[30]), .IN6(
          n737), .Q(n714));
   AO222X1 U970 (.IN1(n501), .IN2(n511), .IN3(n3), .IN4(n738), .IN5(n739), .IN6(n17), .Q(
          n737));
   NAND4X0 U971 (.IN1(n690), .IN2(n564), .IN3(n740), .IN4(n741), .QN(n739));
   OA222X1 U972 (.IN1(n123), .IN2(n138), .IN3(n658), .IN4(n125), .IN5(n115), .IN6(n146), .
          Q(n741));
   AO21X1 U973 (.IN1(n129), .IN2(n130), .IN3(n548), .Q(n740));
   NAND4X0 U974 (.IN1(n731), .IN2(n711), .IN3(n742), .IN4(n743), .QN(n738));
   OA221X1 U975 (.IN1(n655), .IN2(n118), .IN3(n135), .IN4(n122), .IN5(n744), .Q(n743));
   NAND4X0 U976 (.IN1(n642), .IN2(n565), .IN3(n745), .IN4(n746), .QN(n736));
   OA222X1 U977 (.IN1(n554), .IN2(n135), .IN3(n747), .IN4(n122), .IN5(n522), .IN6(n132), .
          Q(n746));
   NAND4X0 U978 (.IN1(n111), .IN2(n694), .IN3(n678), .IN4(n748), .QN(n735));
   OA22X1 U979 (.IN1(n548), .IN2(n645), .IN3(n123), .IN4(n140), .Q(n748));
   AO222X1 U980 (.IN1(n750), .IN2(n751), .IN3(n752), .IN4(n753), .IN5(n754), .IN6(n170), .
          Q(new_sboxw[26]));
   AO222X1 U981 (.IN1(n528), .IN2(n755), .IN3(n530), .IN4(n756), .IN5(sboxw[30]), .IN6(
          n757), .Q(n754));
   NAND4X0 U982 (.IN1(n541), .IN2(n576), .IN3(n758), .IN4(n759), .QN(n757));
   OA22X1 U983 (.IN1(n3), .IN2(n760), .IN3(n138), .IN4(n126), .Q(n759));
   AO222X1 U984 (.IN1(n508), .IN2(n511), .IN3(n730), .IN4(n125), .IN5(sboxw[27]), .IN6(
          n115), .Q(n762));
   AO221X1 U985 (.IN1(n549), .IN2(n539), .IN3(n667), .IN4(n12), .IN5(n525), .Q(n761));
   NAND3X0 U986 (.IN1(n124), .IN2(n583), .IN3(n572), .QN(n763));
   NAND4X0 U987 (.IN1(n711), .IN2(n764), .IN3(n765), .IN4(n766), .QN(n756));
   OAI21X1 U988 (.IN1(n128), .IN2(n554), .IN3(n663), .QN(n512));
   OR2X1 U989 (.IN1(n119), .IN2(n645), .Q(n765));
   NAND4X0 U990 (.IN1(n702), .IN2(n712), .IN3(n768), .IN4(n769), .QN(n755));
   OA221X1 U991 (.IN1(n140), .IN2(n115), .IN3(n539), .IN4(n130), .IN5(n518), .Q(n769));
   OA22X1 U992 (.IN1(n134), .IN2(n122), .IN3(n12), .IN4(n133), .Q(n768));
   AO22X1 U993 (.IN1(sboxw[29]), .IN2(n771), .IN3(n772), .IN4(n17), .Q(n753));
   AO221X1 U994 (.IN1(n770), .IN2(n118), .IN3(n555), .IN4(n119), .IN5(n773), .Q(n772));
   AO221X1 U995 (.IN1(n774), .IN2(n115), .IN3(n522), .IN4(n525), .IN5(n730), .Q(n773));
   NAND4X0 U996 (.IN1(n666), .IN2(n504), .IN3(n775), .IN4(n776), .QN(n771));
   OA222X1 U997 (.IN1(n120), .IN2(n133), .IN3(n747), .IN4(n123), .IN5(n134), .IN6(n122), .
          Q(n776));
   AND2X1 U998 (.IN1(n113), .IN2(n541), .Q(n775));
   AO22X1 U999 (.IN1(sboxw[29]), .IN2(n778), .IN3(n779), .IN4(n17), .Q(n751));
   NAND4X0 U1000 (.IN1(n544), .IN2(n731), .IN3(n780), .IN4(n781), .QN(n779));
   OA222X1 U1001 (.IN1(n12), .IN2(n140), .IN3(n548), .IN4(n134), .IN5(n141), .IN6(n2), .Q(
          n781));
   AND2X1 U1002 (.IN1(n565), .IN2(n712), .Q(n780));
   NAND4X0 U1003 (.IN1(n642), .IN2(n504), .IN3(n782), .IN4(n783), .QN(n778));
   OA222X1 U1004 (.IN1(n129), .IN2(n2), .IN3(n548), .IN4(n133), .IN5(n539), .IN6(n130), .Q(
          n783));
   AO222X1 U1005 (.IN1(n750), .IN2(n784), .IN3(n752), .IN4(n785), .IN5(n786), .IN6(n170), .
          Q(new_sboxw[25]));
   AO221X1 U1006 (.IN1(n640), .IN2(n787), .IN3(n638), .IN4(n788), .IN5(n789), .Q(n786));
   AO22X1 U1007 (.IN1(n528), .IN2(n790), .IN3(n530), .IN4(n791), .Q(n789));
   OA221X1 U1008 (.IN1(n554), .IN2(n132), .IN3(n120), .IN4(n144), .IN5(n745), .Q(n793));
   OA222X1 U1009 (.IN1(n149), .IN2(n115), .IN3(n118), .IN4(n145), .IN5(n11), .IN6(n129), .
          Q(n792));
   NAND4X0 U1010 (.IN1(n576), .IN2(n130), .IN3(n794), .IN4(n795), .QN(n790));
   OA222X1 U1011 (.IN1(n548), .IN2(n128), .IN3(n118), .IN4(n127), .IN5(n539), .IN6(n134), .
          Q(n795));
   NAND4X0 U1012 (.IN1(n505), .IN2(n130), .IN3(n796), .IN4(n797), .QN(n788));
   OA222X1 U1013 (.IN1(sboxw[27]), .IN2(n2), .IN3(n651), .IN4(n120), .IN5(n539), .IN6(n136)
          , .Q(n797));
   NAND4X0 U1014 (.IN1(n572), .IN2(n764), .IN3(n579), .IN4(n798), .QN(n787));
   OA222X1 U1015 (.IN1(n548), .IN2(n129), .IN3(n138), .IN4(n119), .IN5(n115), .IN6(n130), .
          Q(n798));
   AO222X1 U1016 (.IN1(n734), .IN2(n501), .IN3(n3), .IN4(n799), .IN5(n800), .IN6(n17), .Q(
          n785));
   NAND4X0 U1017 (.IN1(n703), .IN2(n542), .IN3(n801), .IN4(n802), .QN(n800));
   OA221X1 U1018 (.IN1(n11), .IN2(n655), .IN3(n141), .IN4(n119), .IN5(n744), .Q(n802));
   NAND4X0 U1019 (.IN1(n121), .IN2(n124), .IN3(n803), .IN4(n804), .QN(n799));
   OA22X1 U1020 (.IN1(n548), .IN2(n146), .IN3(n522), .IN4(n655), .Q(n804));
   AO221X1 U1021 (.IN1(n3), .IN2(n806), .IN3(n550), .IN4(n501), .IN5(n807), .Q(n784));
   AO21X1 U1022 (.IN1(n808), .IN2(n17), .IN3(n777), .Q(n807));
   NAND3X0 U1023 (.IN1(n712), .IN2(n514), .IN3(n809), .QN(n808));
   OA22X1 U1024 (.IN1(n597), .IN2(n122), .IN3(n509), .IN4(n119), .Q(n809));
   AO221X1 U1025 (.IN1(n770), .IN2(n119), .IN3(n538), .IN4(n122), .IN5(n810), .Q(n806));
   AO21X1 U1026 (.IN1(n522), .IN2(n500), .IN3(n734), .Q(n810));
   AO222X1 U1027 (.IN1(n750), .IN2(n811), .IN3(n752), .IN4(n812), .IN5(n813), .IN6(n170), .
          Q(new_sboxw[24]));
   AO222X1 U1028 (.IN1(n528), .IN2(n814), .IN3(n530), .IN4(n815), .IN5(sboxw[30]), .IN6(
          n816), .Q(n813));
   AO221X1 U1029 (.IN1(n817), .IN2(n17), .IN3(n3), .IN4(n818), .IN5(n749), .Q(n816));
   NAND4X0 U1030 (.IN1(n506), .IN2(n129), .IN3(n819), .IN4(n820), .QN(n818));
   OA222X1 U1031 (.IN1(n655), .IN2(n119), .IN3(n522), .IN4(n145), .IN5(n148), .IN6(n122), .
          Q(n820));
   AO22X1 U1032 (.IN1(n555), .IN2(n125), .IN3(n730), .IN4(n115), .Q(n817));
   NAND4X0 U1033 (.IN1(n510), .IN2(n821), .IN3(n822), .IN4(n694), .QN(n815));
   OR2X1 U1034 (.IN1(n148), .IN2(n517), .Q(n821));
   OA22X1 U1035 (.IN1(n139), .IN2(n125), .IN3(n118), .IN4(sboxw[26]), .Q(n517));
   OA221X1 U1036 (.IN1(n136), .IN2(n118), .IN3(n145), .IN4(n120), .IN5(n133), .Q(n510));
   NAND4X0 U1037 (.IN1(n542), .IN2(n582), .IN3(n823), .IN4(n824), .QN(n814));
   OA221X1 U1038 (.IN1(n508), .IN2(n149), .IN3(n11), .IN4(n146), .IN5(n710), .Q(n824));
   OR2X1 U1039 (.IN1(n2), .IN2(n648), .Q(n823));
   NAND3X0 U1040 (.IN1(n767), .IN2(n825), .IN3(n826), .QN(n812));
   OA222X1 U1041 (.IN1(n128), .IN2(n126), .IN3(sboxw[29]), .IN4(n827), .IN5(n828), .IN6(
          n17), .Q(n826));
   OA221X1 U1042 (.IN1(n522), .IN2(n148), .IN3(n118), .IN4(n145), .IN5(n829), .Q(n828));
   OA221X1 U1043 (.IN1(n539), .IN2(n140), .IN3(n508), .IN4(n145), .IN5(n830), .Q(n827));
   AND2X1 U1044 (.IN1(n130), .IN2(n545), .Q(n830));
   OA22X1 U1045 (.IN1(n130), .IN2(n2), .IN3(n134), .IN4(n115), .Q(n767));
   AO221X1 U1046 (.IN1(n831), .IN2(n17), .IN3(n3), .IN4(n832), .IN5(n833), .Q(n811));
   AO22X1 U1047 (.IN1(n724), .IN2(n501), .IN3(n525), .IN4(n122), .Q(n833));
   NAND4X0 U1048 (.IN1(n678), .IN2(n134), .IN3(n834), .IN4(n835), .QN(n832));
   OA22X1 U1049 (.IN1(n508), .IN2(n146), .IN3(n125), .IN4(n140), .Q(n835));
   AO221X1 U1050 (.IN1(n508), .IN2(n523), .IN3(n511), .IN4(n123), .IN5(n836), .Q(n831));
   AO21X1 U1051 (.IN1(n837), .IN2(n122), .IN3(n805), .Q(n836));
   AO22X1 U1052 (.IN1(n838), .IN2(n110), .IN3(sboxw[23]), .IN4(n839), .Q(new_sboxw[23]));
   AO22X1 U1053 (.IN1(n840), .IN2(n109), .IN3(sboxw[22]), .IN4(n841), .Q(n839));
   AO222X1 U1054 (.IN1(n842), .IN2(n843), .IN3(n15), .IN4(n844), .IN5(n845), .IN6(n16), .Q(
          n841));
   NAND4X0 U1055 (.IN1(n846), .IN2(n847), .IN3(n848), .IN4(n849), .QN(n845));
   AO221X1 U1056 (.IN1(n87), .IN2(n76), .IN3(n853), .IN4(n74), .IN5(n854), .Q(n844));
   NAND4X0 U1057 (.IN1(n855), .IN2(n856), .IN3(n857), .IN4(n858), .QN(n840));
   OA221X1 U1058 (.IN1(n859), .IN2(n104), .IN3(n82), .IN4(n86), .IN5(n860), .Q(n858));
   NAND4X0 U1059 (.IN1(n77), .IN2(n84), .IN3(n862), .IN4(n863), .QN(n861));
   OA22X1 U1060 (.IN1(n10), .IN2(n97), .IN3(n864), .IN4(n86), .Q(n863));
   AO221X1 U1061 (.IN1(n867), .IN2(n9), .IN3(n868), .IN4(n76), .IN5(n869), .Q(n866));
   AO222X1 U1062 (.IN1(n870), .IN2(n871), .IN3(n872), .IN4(n873), .IN5(sboxw[22]), .IN6(
          n874), .Q(n838));
   AO221X1 U1063 (.IN1(n875), .IN2(n16), .IN3(n865), .IN4(n843), .IN5(n876), .Q(n874));
   AO21X1 U1064 (.IN1(n15), .IN2(n877), .IN3(n878), .Q(n876));
   AO221X1 U1065 (.IN1(n879), .IN2(n71), .IN3(n880), .IN4(n881), .IN5(n882), .Q(n877));
   NAND4X0 U1066 (.IN1(n883), .IN2(n92), .IN3(n884), .IN4(n885), .QN(n875));
   OA22X1 U1067 (.IN1(n9), .IN2(n83), .IN3(n850), .IN4(n96), .Q(n885));
   NAND4X0 U1068 (.IN1(n886), .IN2(n887), .IN3(n888), .IN4(n889), .QN(n873));
   OA22X1 U1069 (.IN1(n10), .IN2(n94), .IN3(n850), .IN4(n91), .Q(n889));
   AO221X1 U1070 (.IN1(n890), .IN2(n891), .IN3(n892), .IN4(n864), .IN5(n893), .Q(n871));
   AO221X1 U1071 (.IN1(n894), .IN2(n74), .IN3(n895), .IN4(n896), .IN5(n897), .Q(n893));
   AO222X1 U1072 (.IN1(n898), .IN2(n899), .IN3(n900), .IN4(n901), .IN5(sboxw[23]), .IN6(
          n902), .Q(new_sboxw[22]));
   AO222X1 U1073 (.IN1(n872), .IN2(n903), .IN3(sboxw[22]), .IN4(n904), .IN5(n870), .IN6(
          n905), .Q(n902));
   NAND4X0 U1074 (.IN1(n906), .IN2(n907), .IN3(n908), .IN4(n909), .QN(n905));
   OA221X1 U1075 (.IN1(n104), .IN2(n71), .IN3(n97), .IN4(n78), .IN5(n910), .Q(n909));
   OA22X1 U1076 (.IN1(n79), .IN2(n83), .IN3(n890), .IN4(n88), .Q(n908));
   NAND4X0 U1078 (.IN1(n913), .IN2(n914), .IN3(n915), .IN4(n916), .QN(n912));
   OA222X1 U1079 (.IN1(n917), .IN2(n105), .IN3(n76), .IN4(n89), .IN5(n84), .IN6(n71), .Q(
          n916));
   AND2X1 U1080 (.IN1(n918), .IN2(n919), .Q(n915));
   NAND4X0 U1081 (.IN1(n920), .IN2(n921), .IN3(n922), .IN4(n923), .QN(n911));
   AND4X1 U1082 (.IN1(n907), .IN2(n924), .IN3(n925), .IN4(n919), .Q(n923));
   OA22X1 U1083 (.IN1(n74), .IN2(n102), .IN3(n10), .IN4(n84), .Q(n922));
   NAND4X0 U1084 (.IN1(n919), .IN2(n887), .IN3(n927), .IN4(n928), .QN(n903));
   OA22X1 U1085 (.IN1(n896), .IN2(n92), .IN3(n881), .IN4(n101), .Q(n928));
   NAND4X0 U1087 (.IN1(n856), .IN2(n89), .IN3(n931), .IN4(n932), .QN(n930));
   OA222X1 U1088 (.IN1(n881), .IN2(n91), .IN3(n10), .IN4(n97), .IN5(n890), .IN6(n96), .Q(
          n932));
   OA22X1 U1089 (.IN1(n92), .IN2(n78), .IN3(n81), .IN4(n101), .Q(n931));
   NAND4X0 U1090 (.IN1(n907), .IN2(n90), .IN3(n70), .IN4(n933), .QN(n929));
   OA222X1 U1091 (.IN1(n9), .IN2(n91), .IN3(n10), .IN4(n99), .IN5(n74), .IN6(n83), .Q(n933)
          );
   NAND3X0 U1092 (.IN1(n913), .IN2(n934), .IN3(n935), .QN(n899));
   OA22X1 U1093 (.IN1(n936), .IN2(n16), .IN3(n15), .IN4(n937), .Q(n935));
   OA221X1 U1094 (.IN1(n104), .IN2(n74), .IN3(n10), .IN4(n90), .IN5(n938), .Q(n937));
   OA22X1 U1095 (.IN1(n864), .IN2(n105), .IN3(sboxw[18]), .IN4(n890), .Q(n938));
   OA221X1 U1096 (.IN1(n917), .IN2(n102), .IN3(n939), .IN4(n79), .IN5(n919), .Q(n936));
   AO222X1 U1097 (.IN1(n898), .IN2(n940), .IN3(n900), .IN4(n941), .IN5(sboxw[23]), .IN6(
          n942), .Q(new_sboxw[21]));
   AO221X1 U1098 (.IN1(n872), .IN2(n943), .IN3(n870), .IN4(n944), .IN5(n945), .Q(n942));
   AO22X1 U1099 (.IN1(n946), .IN2(n947), .IN3(n948), .IN4(n949), .Q(n945));
   NAND4X0 U1100 (.IN1(n950), .IN2(n847), .IN3(n951), .IN4(n952), .QN(n949));
   OA222X1 U1101 (.IN1(n896), .IN2(n85), .IN3(n74), .IN4(n86), .IN5(n81), .IN6(n96), .Q(
          n952));
   OA22X1 U1102 (.IN1(n953), .IN2(n71), .IN3(n9), .IN4(n90), .Q(n951));
   NAND3X0 U1103 (.IN1(n910), .IN2(n954), .IN3(n955), .QN(n947));
   OA221X1 U1104 (.IN1(n896), .IN2(n104), .IN3(n10), .IN4(n956), .IN5(n957), .Q(n955));
   NAND3X0 U1105 (.IN1(n958), .IN2(n959), .IN3(n960), .QN(n944));
   OA221X1 U1106 (.IN1(n881), .IN2(n98), .IN3(n961), .IN4(n76), .IN5(n962), .Q(n960));
   OA22X1 U1107 (.IN1(n79), .IN2(n96), .IN3(n963), .IN4(n74), .Q(n958));
   NAND4X0 U1108 (.IN1(n69), .IN2(n924), .IN3(n964), .IN4(n965), .QN(n943));
   OA222X1 U1109 (.IN1(n896), .IN2(n84), .IN3(n94), .IN4(n74), .IN5(n81), .IN6(n86), .Q(
          n965));
   NAND4X0 U1111 (.IN1(n970), .IN2(n971), .IN3(n972), .IN4(n973), .QN(n969));
   AND4X1 U1112 (.IN1(n94), .IN2(n887), .IN3(n77), .IN4(n974), .Q(n973));
   OA22X1 U1113 (.IN1(n850), .IN2(n83), .IN3(n76), .IN4(n88), .Q(n972));
   NAND4X0 U1114 (.IN1(n967), .IN2(n80), .IN3(n976), .IN4(n977), .QN(n968));
   OA222X1 U1115 (.IN1(n9), .IN2(n85), .IN3(n890), .IN4(n83), .IN5(n74), .IN6(n90), .Q(
          n977));
   AND2X1 U1116 (.IN1(n924), .IN2(n847), .Q(n976));
   AO221X1 U1117 (.IN1(n865), .IN2(n843), .IN3(n978), .IN4(n73), .IN5(n979), .Q(n940));
   AO221X1 U1118 (.IN1(n15), .IN2(n980), .IN3(n981), .IN4(n16), .IN5(n72), .Q(n979));
   NAND3X0 U1119 (.IN1(n896), .IN2(n15), .IN3(n982), .QN(n934));
   NAND4X0 U1120 (.IN1(n921), .IN2(n96), .IN3(n983), .IN4(n984), .QN(n981));
   AO222X1 U1121 (.IN1(n898), .IN2(n988), .IN3(n900), .IN4(n989), .IN5(sboxw[23]), .IN6(
          n990), .Q(new_sboxw[20]));
   AO221X1 U1122 (.IN1(n948), .IN2(n991), .IN3(n946), .IN4(n992), .IN5(n993), .Q(n990));
   AO22X1 U1123 (.IN1(n870), .IN2(n994), .IN3(n872), .IN4(n995), .Q(n993));
   NAND4X0 U1124 (.IN1(n856), .IN2(n925), .IN3(n974), .IN4(n996), .QN(n995));
   AOI222X1 U1125 (.IN1(n881), .IN2(n853), .IN3(n79), .IN4(n997), .IN5(n867), .IN6(n987), .
          QN(n996));
   NAND4X0 U1126 (.IN1(n998), .IN2(n918), .IN3(n999), .IN4(n1000), .QN(n994));
   OA222X1 U1127 (.IN1(n10), .IN2(n84), .IN3(n864), .IN4(n90), .IN5(n896), .IN6(n89), .Q(
          n1000));
   NAND4X0 U1128 (.IN1(n967), .IN2(n1002), .IN3(n1003), .IN4(n1004), .QN(n992));
   OA221X1 U1129 (.IN1(n81), .IN2(n94), .IN3(n97), .IN4(n75), .IN5(n985), .Q(n1004));
   AO21X1 U1130 (.IN1(n85), .IN2(n96), .IN3(n78), .Q(n1003));
   OA221X1 U1131 (.IN1(n850), .IN2(n97), .IN3(n864), .IN4(n99), .IN5(n957), .Q(n1006));
   OA222X1 U1132 (.IN1(n963), .IN2(n81), .IN3(n9), .IN4(n89), .IN5(n10), .IN6(n86), .Q(
          n1005));
   AO222X1 U1133 (.IN1(n1007), .IN2(n16), .IN3(n15), .IN4(n1008), .IN5(n843), .IN6(n869), .
          Q(n989));
   NAND4X0 U1134 (.IN1(n77), .IN2(n96), .IN3(n886), .IN4(n1009), .QN(n1008));
   OA22X1 U1135 (.IN1(n987), .IN2(n102), .IN3(n94), .IN4(n71), .Q(n1009));
   NAND4X0 U1136 (.IN1(n1010), .IN2(n1011), .IN3(n1012), .IN4(n1013), .QN(n1007));
   OA222X1 U1137 (.IN1(n9), .IN2(n105), .IN3(n74), .IN4(n89), .IN5(n96), .IN6(n75), .Q(
          n1013));
   AO222X1 U1138 (.IN1(n843), .IN2(n997), .IN3(n15), .IN4(n1014), .IN5(n1015), .IN6(n16), .
          Q(n988));
   NAND4X0 U1139 (.IN1(n77), .IN2(n998), .IN3(n1016), .IN4(n1017), .QN(n1015));
   OA221X1 U1140 (.IN1(n81), .IN2(n94), .IN3(n890), .IN4(n1018), .IN5(n1019), .Q(n1017));
   AND2X1 U1141 (.IN1(n907), .IN2(n887), .Q(n1016));
   NAND4X0 U1142 (.IN1(n1020), .IN2(n887), .IN3(n1001), .IN4(n1021), .QN(n1014));
   OA22X1 U1143 (.IN1(n987), .IN2(n101), .IN3(n74), .IN4(n86), .Q(n1021));
   OA22X1 U1144 (.IN1(n78), .IN2(sboxw[18]), .IN3(n74), .IN4(n95), .Q(n987));
   AO222X1 U1145 (.IN1(n598), .IN2(n1022), .IN3(n600), .IN4(n1023), .IN5(n1024), .IN6(
          n1408), .Q(new_sboxw[1]));
   AO221X1 U1146 (.IN1(n386), .IN2(n1025), .IN3(n384), .IN4(n1026), .IN5(n1027), .Q(n1024)
          );
   AO22X1 U1147 (.IN1(n308), .IN2(n1028), .IN3(n310), .IN4(n1029), .Q(n1027));
   OA221X1 U1148 (.IN1(n334), .IN2(n156), .IN3(n27), .IN4(n168), .IN5(n491), .Q(n1031));
   OA222X1 U1149 (.IN1(n1405), .IN2(n22), .IN3(n25), .IN4(n171), .IN5(n4), .IN6(n153), .Q(
          n1030));
   NAND4X0 U1150 (.IN1(n356), .IN2(n154), .IN3(n1032), .IN4(n1033), .QN(n1028));
   OA222X1 U1151 (.IN1(n328), .IN2(n152), .IN3(n25), .IN4(n151), .IN5(n319), .IN6(n158), .
          Q(n1033));
   NAND4X0 U1152 (.IN1(n285), .IN2(n154), .IN3(n1034), .IN4(n1035), .QN(n1026));
   OA222X1 U1153 (.IN1(sboxw[3]), .IN2(n29), .IN3(n397), .IN4(n27), .IN5(n319), .IN6(n160)
          , .Q(n1035));
   NAND4X0 U1154 (.IN1(n352), .IN2(n612), .IN3(n359), .IN4(n1036), .QN(n1025));
   OA222X1 U1155 (.IN1(n328), .IN2(n153), .IN3(n162), .IN4(n26), .IN5(n22), .IN6(n154), .Q(
          n1036));
   AO222X1 U1156 (.IN1(n480), .IN2(n281), .IN3(n13), .IN4(n1037), .IN5(n1038), .IN6(n14), .
          Q(n1023));
   NAND4X0 U1157 (.IN1(n449), .IN2(n322), .IN3(n1039), .IN4(n1040), .QN(n1038));
   OA221X1 U1158 (.IN1(n4), .IN2(n401), .IN3(n165), .IN4(n26), .IN5(n490), .Q(n1040));
   NAND4X0 U1159 (.IN1(n28), .IN2(n31), .IN3(n1041), .IN4(n1042), .QN(n1037));
   OA22X1 U1160 (.IN1(n328), .IN2(n1402), .IN3(n302), .IN4(n401), .Q(n1042));
   AO221X1 U1161 (.IN1(n13), .IN2(n1044), .IN3(n330), .IN4(n281), .IN5(n1045), .Q(n1022)
          );
   AO21X1 U1162 (.IN1(n1046), .IN2(n14), .IN3(n625), .Q(n1045));
   NAND3X0 U1163 (.IN1(n458), .IN2(n294), .IN3(n1047), .QN(n1046));
   OA22X1 U1164 (.IN1(n377), .IN2(n29), .IN3(n289), .IN4(n26), .Q(n1047));
   AO221X1 U1165 (.IN1(n618), .IN2(n26), .IN3(n318), .IN4(n29), .IN5(n1048), .Q(n1044));
   AO21X1 U1166 (.IN1(n302), .IN2(n280), .IN3(n480), .Q(n1048));
   AO22X1 U1167 (.IN1(sboxw[23]), .IN2(n1049), .IN3(n1050), .IN4(n110), .Q(new_sboxw[19])
          );
   AO222X1 U1168 (.IN1(n946), .IN2(n1051), .IN3(n948), .IN4(n1052), .IN5(n1053), .IN6(n109)
          , .Q(n1050));
   AO222X1 U1169 (.IN1(n843), .IN2(n93), .IN3(n15), .IN4(n1054), .IN5(n1055), .IN6(n16), .
          Q(n1053));
   NAND4X0 U1170 (.IN1(n1056), .IN2(n1001), .IN3(n1057), .IN4(n1058), .QN(n1055));
   AND3X1 U1171 (.IN1(n906), .IN2(n957), .IN3(n1010), .Q(n1058));
   NAND4X0 U1172 (.IN1(n1060), .IN2(n883), .IN3(n67), .IN4(n957), .QN(n1054));
   OR2X1 U1173 (.IN1(n74), .IN2(n851), .Q(n1060));
   NAND4X0 U1174 (.IN1(n1002), .IN2(n86), .IN3(n913), .IN4(n1062), .QN(n1052));
   OA222X1 U1175 (.IN1(n9), .IN2(n105), .IN3(n850), .IN4(n1063), .IN5(n959), .IN6(n79), .Q(
          n1062));
   NAND4X0 U1176 (.IN1(n1066), .IN2(n1011), .IN3(n1067), .IN4(n1068), .QN(n1051));
   OA221X1 U1177 (.IN1(n84), .IN2(n78), .IN3(n79), .IN4(n90), .IN5(n1057), .Q(n1068));
   AND2X1 U1178 (.IN1(n918), .IN2(n80), .Q(n1067));
   AO222X1 U1179 (.IN1(n870), .IN2(n1070), .IN3(n872), .IN4(n1071), .IN5(sboxw[22]), .IN6(
          n1072), .Q(n1049));
   AO222X1 U1180 (.IN1(n843), .IN2(n853), .IN3(n15), .IN4(n1073), .IN5(n1074), .IN6(n16), .
          Q(n1072));
   NAND4X0 U1181 (.IN1(n998), .IN2(n906), .IN3(n1075), .IN4(n1076), .QN(n1074));
   OA222X1 U1182 (.IN1(n79), .IN2(n94), .IN3(n966), .IN4(n81), .IN5(n71), .IN6(n102), .Q(
          n1076));
   AO21X1 U1183 (.IN1(n85), .IN2(n86), .IN3(n890), .Q(n1075));
   NAND4X0 U1184 (.IN1(n1066), .IN2(n1019), .IN3(n1077), .IN4(n1078), .QN(n1073));
   OA221X1 U1185 (.IN1(n963), .IN2(n74), .IN3(n91), .IN4(n78), .IN5(n1079), .Q(n1078));
   NAND4X0 U1186 (.IN1(n950), .IN2(n907), .IN3(n1080), .IN4(n1081), .QN(n1071));
   OA222X1 U1187 (.IN1(n896), .IN2(n91), .IN3(n1082), .IN4(n78), .IN5(n864), .IN6(n88), .Q(
          n1081));
   NAND4X0 U1188 (.IN1(n67), .IN2(n1002), .IN3(n986), .IN4(n1083), .QN(n1070));
   OA22X1 U1189 (.IN1(n890), .IN2(n953), .IN3(n79), .IN4(n96), .Q(n1083));
   AO222X1 U1190 (.IN1(n1085), .IN2(n1086), .IN3(n1087), .IN4(n1088), .IN5(n1089), .IN6(
          n110), .Q(new_sboxw[18]));
   AO222X1 U1191 (.IN1(n870), .IN2(n1090), .IN3(n872), .IN4(n1091), .IN5(sboxw[22]), .IN6(
          n1092), .Q(n1089));
   NAND4X0 U1192 (.IN1(n883), .IN2(n918), .IN3(n1093), .IN4(n1094), .QN(n1092));
   OA22X1 U1193 (.IN1(n15), .IN2(n1095), .IN3(n94), .IN4(n82), .Q(n1094));
   AO222X1 U1194 (.IN1(n850), .IN2(n853), .IN3(n1065), .IN4(n81), .IN5(sboxw[19]), .IN6(
          n71), .Q(n1097));
   AO221X1 U1195 (.IN1(n891), .IN2(n881), .IN3(n975), .IN4(n10), .IN5(n867), .Q(n1096));
   NAND3X0 U1196 (.IN1(n80), .IN2(n925), .IN3(n914), .QN(n1098));
   NAND4X0 U1197 (.IN1(n1019), .IN2(n1099), .IN3(n1100), .IN4(n1101), .QN(n1091));
   OAI21X1 U1198 (.IN1(n84), .IN2(n896), .IN3(n971), .QN(n854));
   OR2X1 U1199 (.IN1(n75), .IN2(n953), .Q(n1100));
   NAND4X0 U1200 (.IN1(n1010), .IN2(n1020), .IN3(n1103), .IN4(n1104), .QN(n1090));
   OA221X1 U1201 (.IN1(n96), .IN2(n71), .IN3(n881), .IN4(n86), .IN5(n860), .Q(n1104));
   OA22X1 U1202 (.IN1(n90), .IN2(n78), .IN3(n10), .IN4(n89), .Q(n1103));
   AO221X1 U1204 (.IN1(n1105), .IN2(n74), .IN3(n897), .IN4(n75), .IN5(n1108), .Q(n1107));
   AO221X1 U1205 (.IN1(n1109), .IN2(n71), .IN3(n864), .IN4(n867), .IN5(n1065), .Q(n1108)
          );
   NAND4X0 U1206 (.IN1(n974), .IN2(n846), .IN3(n1110), .IN4(n1111), .QN(n1106));
   OA222X1 U1207 (.IN1(n76), .IN2(n89), .IN3(n1082), .IN4(n79), .IN5(n90), .IN6(n78), .Q(
          n1111));
   AND2X1 U1208 (.IN1(n69), .IN2(n883), .Q(n1110));
   NAND4X0 U1210 (.IN1(n886), .IN2(n1066), .IN3(n1115), .IN4(n1116), .QN(n1114));
   OA222X1 U1211 (.IN1(n10), .IN2(n96), .IN3(n890), .IN4(n90), .IN5(n97), .IN6(n78), .Q(
          n1116));
   AND2X1 U1212 (.IN1(n907), .IN2(n1020), .Q(n1115));
   NAND4X0 U1213 (.IN1(n950), .IN2(n846), .IN3(n1117), .IN4(n1118), .QN(n1113));
   OA222X1 U1214 (.IN1(n85), .IN2(n78), .IN3(n890), .IN4(n89), .IN5(n881), .IN6(n86), .Q(
          n1118));
   AO222X1 U1215 (.IN1(n1085), .IN2(n1119), .IN3(n1087), .IN4(n1120), .IN5(n1121), .IN6(
          n110), .Q(new_sboxw[17]));
   AO221X1 U1216 (.IN1(n948), .IN2(n1122), .IN3(n946), .IN4(n1123), .IN5(n1124), .Q(n1121)
          );
   AO22X1 U1217 (.IN1(n870), .IN2(n1125), .IN3(n872), .IN4(n1126), .Q(n1124));
   OA221X1 U1218 (.IN1(n896), .IN2(n88), .IN3(n76), .IN4(n100), .IN5(n1080), .Q(n1128));
   OA222X1 U1219 (.IN1(n105), .IN2(n71), .IN3(n74), .IN4(n101), .IN5(n9), .IN6(n85), .Q(
          n1127));
   NAND4X0 U1220 (.IN1(n918), .IN2(n86), .IN3(n1129), .IN4(n1130), .QN(n1125));
   OA222X1 U1221 (.IN1(n890), .IN2(n84), .IN3(n74), .IN4(n83), .IN5(n881), .IN6(n90), .Q(
          n1130));
   NAND4X0 U1222 (.IN1(n847), .IN2(n86), .IN3(n1131), .IN4(n1132), .QN(n1123));
   OA222X1 U1223 (.IN1(sboxw[19]), .IN2(n78), .IN3(n959), .IN4(n76), .IN5(n881), .IN6(n92)
          , .Q(n1132));
   NAND4X0 U1224 (.IN1(n914), .IN2(n1099), .IN3(n921), .IN4(n1133), .QN(n1122));
   OA222X1 U1225 (.IN1(n890), .IN2(n85), .IN3(n94), .IN4(n75), .IN5(n71), .IN6(n86), .Q(
          n1133));
   AO222X1 U1226 (.IN1(n1069), .IN2(n843), .IN3(n15), .IN4(n1134), .IN5(n1135), .IN6(n16)
          , .Q(n1120));
   NAND4X0 U1227 (.IN1(n1011), .IN2(n884), .IN3(n1136), .IN4(n1137), .QN(n1135));
   OA221X1 U1228 (.IN1(n9), .IN2(n963), .IN3(n97), .IN4(n75), .IN5(n1079), .Q(n1137));
   NAND4X0 U1229 (.IN1(n77), .IN2(n80), .IN3(n1138), .IN4(n1139), .QN(n1134));
   OA22X1 U1230 (.IN1(n890), .IN2(n102), .IN3(n864), .IN4(n963), .Q(n1139));
   AO221X1 U1231 (.IN1(n15), .IN2(n1141), .IN3(n892), .IN4(n843), .IN5(n1142), .Q(n1119)
          );
   AO21X1 U1232 (.IN1(n1143), .IN2(n16), .IN3(n1112), .Q(n1142));
   NAND3X0 U1233 (.IN1(n1020), .IN2(n856), .IN3(n1144), .QN(n1143));
   OA22X1 U1234 (.IN1(n939), .IN2(n78), .IN3(n851), .IN4(n75), .Q(n1144));
   AO221X1 U1235 (.IN1(n1105), .IN2(n75), .IN3(n880), .IN4(n78), .IN5(n1145), .Q(n1141));
   AO21X1 U1236 (.IN1(n864), .IN2(n842), .IN3(n1069), .Q(n1145));
   AO222X1 U1237 (.IN1(n1085), .IN2(n1146), .IN3(n1087), .IN4(n1147), .IN5(n1148), .IN6(
          n110), .Q(new_sboxw[16]));
   AO222X1 U1238 (.IN1(n870), .IN2(n1149), .IN3(n872), .IN4(n1150), .IN5(sboxw[22]), .IN6(
          n1151), .Q(n1148));
   AO221X1 U1239 (.IN1(n1152), .IN2(n16), .IN3(n15), .IN4(n1153), .IN5(n1084), .Q(n1151)
          );
   NAND4X0 U1240 (.IN1(n848), .IN2(n85), .IN3(n1154), .IN4(n1155), .QN(n1153));
   OA222X1 U1241 (.IN1(n963), .IN2(n75), .IN3(n864), .IN4(n101), .IN5(n104), .IN6(n78), .Q(
          n1155));
   AO22X1 U1242 (.IN1(n897), .IN2(n81), .IN3(n1065), .IN4(n71), .Q(n1152));
   NAND4X0 U1243 (.IN1(n852), .IN2(n1156), .IN3(n1157), .IN4(n1002), .QN(n1150));
   OR2X1 U1244 (.IN1(n104), .IN2(n859), .Q(n1156));
   OA22X1 U1245 (.IN1(n95), .IN2(n81), .IN3(n74), .IN4(sboxw[18]), .Q(n859));
   OA221X1 U1246 (.IN1(n92), .IN2(n74), .IN3(n101), .IN4(n76), .IN5(n89), .Q(n852));
   NAND4X0 U1247 (.IN1(n884), .IN2(n924), .IN3(n1158), .IN4(n1159), .QN(n1149));
   OA221X1 U1248 (.IN1(n850), .IN2(n105), .IN3(n9), .IN4(n102), .IN5(n1018), .Q(n1159));
   OR2X1 U1249 (.IN1(n78), .IN2(n956), .Q(n1158));
   NAND3X0 U1250 (.IN1(n1102), .IN2(n1160), .IN3(n1161), .QN(n1147));
   OA221X1 U1252 (.IN1(n864), .IN2(n104), .IN3(n74), .IN4(n101), .IN5(n1164), .Q(n1163));
   OA221X1 U1253 (.IN1(n881), .IN2(n96), .IN3(n850), .IN4(n101), .IN5(n1165), .Q(n1162));
   AND2X1 U1254 (.IN1(n86), .IN2(n887), .Q(n1165));
   OA22X1 U1255 (.IN1(n86), .IN2(n78), .IN3(n90), .IN4(n71), .Q(n1102));
   AO221X1 U1256 (.IN1(n1166), .IN2(n16), .IN3(n15), .IN4(n1167), .IN5(n1168), .Q(n1146)
          );
   AO22X1 U1257 (.IN1(n1059), .IN2(n843), .IN3(n867), .IN4(n78), .Q(n1168));
   NAND4X0 U1258 (.IN1(n986), .IN2(n90), .IN3(n1169), .IN4(n1170), .QN(n1167));
   OA22X1 U1259 (.IN1(n850), .IN2(n102), .IN3(n81), .IN4(n96), .Q(n1170));
   AO221X1 U1260 (.IN1(n850), .IN2(n865), .IN3(n853), .IN4(n79), .IN5(n1171), .Q(n1166));
   AO21X1 U1261 (.IN1(n1172), .IN2(n78), .IN3(n1140), .Q(n1171));
   AO22X1 U1262 (.IN1(n1173), .IN2(n66), .IN3(sboxw[15]), .IN4(n1174), .Q(new_sboxw[15])
          );
   OAI22X1 U1263 (.IN1(sboxw[14]), .IN2(n1175), .IN3(n1176), .IN4(n65), .QN(n1174));
   OA222X1 U1264 (.IN1(n8), .IN2(n1177), .IN3(n1178), .IN4(n64), .IN5(n63), .IN6(n53), .Q(
          n1176));
   OA221X1 U1265 (.IN1(n193), .IN2(n37), .IN3(n6), .IN4(n244), .IN5(n1179), .Q(n1178));
   AND4X1 U1266 (.IN1(n1180), .IN2(n1181), .IN3(n197), .IN4(n1182), .Q(n1177));
   AND3X1 U1267 (.IN1(n241), .IN2(n1183), .IN3(n245), .Q(n1180));
   OA221X1 U1268 (.IN1(n35), .IN2(n1409), .IN3(n58), .IN4(n1412), .IN5(n41), .Q(n245));
   AO221X1 U1269 (.IN1(n205), .IN2(n206), .IN3(n250), .IN4(n251), .IN5(n44), .Q(n1186));
   AO22X1 U1270 (.IN1(n7), .IN2(sboxw[10]), .IN3(n193), .IN4(n48), .Q(n251));
   AO221X1 U1271 (.IN1(n8), .IN2(n1188), .IN3(n1189), .IN4(n64), .IN5(n1190), .Q(n1185));
   NAND4X0 U1272 (.IN1(n40), .IN2(n46), .IN3(n1191), .IN4(n1192), .QN(n1189));
   OA22X1 U1273 (.IN1(n7), .IN2(n51), .IN3(n219), .IN4(n47), .Q(n1192));
   AO221X1 U1274 (.IN1(n269), .IN2(n6), .IN3(n1193), .IN4(n1412), .IN5(n238), .Q(n1188));
   AO222X1 U1275 (.IN1(n182), .IN2(n1194), .IN3(n184), .IN4(n1195), .IN5(sboxw[14]), .IN6(
          n1196), .Q(n1173));
   AO221X1 U1276 (.IN1(n1197), .IN2(n64), .IN3(n206), .IN4(n273), .IN5(n1198), .Q(n1196)
          );
   AO21X1 U1277 (.IN1(n8), .IN2(n1199), .IN3(n1200), .Q(n1198));
   AO221X1 U1278 (.IN1(n1201), .IN2(n1411), .IN3(n194), .IN4(n1202), .IN5(n262), .Q(n1199)
          );
   NAND4X0 U1279 (.IN1(n1203), .IN2(n35), .IN3(n1182), .IN4(n1204), .QN(n1197));
   NAND4X0 U1280 (.IN1(n1205), .IN2(n264), .IN3(n1183), .IN4(n1206), .QN(n1195));
   OA22X1 U1281 (.IN1(sboxw[10]), .IN2(n1414), .IN3(n7), .IN4(n37), .Q(n1206));
   AO221X1 U1282 (.IN1(n1207), .IN2(n188), .IN3(n221), .IN4(n219), .IN5(n1208), .Q(n1194)
          );
   AO221X1 U1283 (.IN1(n1209), .IN2(n1409), .IN3(n1184), .IN4(n193), .IN5(n239), .Q(n1208)
          );
   AO222X1 U1284 (.IN1(n1210), .IN2(n1211), .IN3(n1212), .IN4(n1213), .IN5(sboxw[15]), .
          IN6(n1214), .Q(new_sboxw[14]));
   AO222X1 U1285 (.IN1(n184), .IN2(n1215), .IN3(sboxw[14]), .IN4(n1216), .IN5(n182), .IN6(
          n1217), .Q(n1214));
   NAND4X0 U1286 (.IN1(n1218), .IN2(n1219), .IN3(n1220), .IN4(n1221), .QN(n1217));
   OA221X1 U1287 (.IN1(n61), .IN2(n1411), .IN3(n51), .IN4(n1414), .IN5(n1222), .Q(n1221)
          );
   OA22X1 U1288 (.IN1(n1413), .IN2(n34), .IN3(n193), .IN4(n33), .Q(n1220));
   AO22X1 U1289 (.IN1(n8), .IN2(n1223), .IN3(n1224), .IN4(n64), .Q(n1216));
   NAND4X0 U1290 (.IN1(n202), .IN2(n1225), .IN3(n1226), .IN4(n1227), .QN(n1224));
   OA222X1 U1291 (.IN1(n1228), .IN2(n60), .IN3(n41), .IN4(n1412), .IN5(n1411), .IN6(n46), .
          Q(n1227));
   AND2X1 U1292 (.IN1(n190), .IN2(n52), .Q(n1226));
   NAND4X0 U1293 (.IN1(n203), .IN2(n1225), .IN3(n1229), .IN4(n1230), .QN(n1223));
   OA222X1 U1294 (.IN1(n7), .IN2(n46), .IN3(n249), .IN4(n1411), .IN5(n1231), .IN6(n1412), .
          Q(n1230));
   AND2X1 U1295 (.IN1(n1219), .IN2(n1232), .Q(n1229));
   NAND4X0 U1296 (.IN1(n1225), .IN2(n264), .IN3(n1233), .IN4(n1234), .QN(n1215));
   OA22X1 U1297 (.IN1(n188), .IN2(n35), .IN3(n194), .IN4(n58), .Q(n1234));
   AO22X1 U1298 (.IN1(n8), .IN2(n1235), .IN3(n1236), .IN4(n64), .Q(n1213));
   NAND4X0 U1299 (.IN1(n45), .IN2(n41), .IN3(n1237), .IN4(n1238), .QN(n1236));
   OA222X1 U1300 (.IN1(n194), .IN2(n42), .IN3(n7), .IN4(n51), .IN5(n193), .IN6(n53), .Q(
          n1238));
   OA22X1 U1301 (.IN1(n1), .IN2(n35), .IN3(n1415), .IN4(n58), .Q(n1237));
   NAND4X0 U1302 (.IN1(n1219), .IN2(n38), .IN3(n50), .IN4(n1239), .QN(n1235));
   OA222X1 U1303 (.IN1(n6), .IN2(n42), .IN3(n7), .IN4(n49), .IN5(n1409), .IN6(n34), .Q(
          n1239));
   AO221X1 U1304 (.IN1(n1240), .IN2(n64), .IN3(n8), .IN4(n1241), .IN5(n1242), .Q(n1211));
   NAND4X0 U1305 (.IN1(n54), .IN2(n1225), .IN3(n1243), .IN4(n1244), .QN(n1241));
   OA22X1 U1306 (.IN1(n41), .IN2(n1411), .IN3(n60), .IN4(n1413), .Q(n1244));
   OR2X1 U1307 (.IN1(n57), .IN2(n1228), .Q(n1243));
   AO221X1 U1308 (.IN1(n1202), .IN2(n1), .IN3(n1409), .IN4(n48), .IN5(n1246), .Q(n1240));
   AO22X1 U1309 (.IN1(n193), .IN2(n250), .IN3(n1193), .IN4(n1415), .Q(n1246));
   AO222X1 U1310 (.IN1(n1210), .IN2(n1247), .IN3(n1212), .IN4(n1248), .IN5(sboxw[15]), .
          IN6(n1249), .Q(new_sboxw[13]));
   AO221X1 U1311 (.IN1(n184), .IN2(n1250), .IN3(n182), .IN4(n1251), .IN5(n1252), .Q(n1249)
          );
   AO22X1 U1312 (.IN1(n179), .IN2(n1253), .IN3(n177), .IN4(n1254), .Q(n1252));
   NAND4X0 U1313 (.IN1(n1255), .IN2(n197), .IN3(n1256), .IN4(n1257), .QN(n1254));
   OA222X1 U1314 (.IN1(n188), .IN2(n43), .IN3(n47), .IN4(n1409), .IN5(n1415), .IN6(n53), .
          Q(n1257));
   OA22X1 U1315 (.IN1(n193), .IN2(n51), .IN3(n6), .IN4(n38), .Q(n1256));
   NAND3X0 U1316 (.IN1(n1222), .IN2(n1259), .IN3(n1260), .QN(n1253));
   OA221X1 U1317 (.IN1(n188), .IN2(n61), .IN3(n7), .IN4(n254), .IN5(n1261), .Q(n1260));
   NAND3X0 U1318 (.IN1(n1263), .IN2(n200), .IN3(n1264), .QN(n1251));
   OA221X1 U1319 (.IN1(n194), .IN2(n55), .IN3(n1265), .IN4(n1412), .IN5(n1266), .Q(n1264)
          );
   OA22X1 U1320 (.IN1(n1413), .IN2(n53), .IN3(n213), .IN4(n1409), .Q(n1263));
   NAND3X0 U1321 (.IN1(n1267), .IN2(n1268), .IN3(n1269), .QN(n1250));
   OA221X1 U1322 (.IN1(n37), .IN2(n1409), .IN3(n6), .IN4(n1270), .IN5(n224), .Q(n1269));
   OA22X1 U1323 (.IN1(n1415), .IN2(n47), .IN3(n188), .IN4(n46), .Q(n1267));
   AO22X1 U1324 (.IN1(n8), .IN2(n1271), .IN3(n1272), .IN4(n64), .Q(n1248));
   NAND4X0 U1325 (.IN1(n1273), .IN2(n1274), .IN3(n1275), .IN4(n1276), .QN(n1272));
   AND4X1 U1326 (.IN1(n37), .IN2(n264), .IN3(n40), .IN4(n1277), .Q(n1276));
   OA22X1 U1327 (.IN1(n225), .IN2(n34), .IN3(n1412), .IN4(n33), .Q(n1275));
   NAND4X0 U1328 (.IN1(n216), .IN2(n197), .IN3(n1278), .IN4(n1279), .QN(n1271));
   OA221X1 U1329 (.IN1(n6), .IN2(n43), .IN3(n1409), .IN4(n38), .IN5(n1268), .Q(n1279));
   OA22X1 U1330 (.IN1(n53), .IN2(n1412), .IN3(n1410), .IN4(n41), .Q(n1268));
   AO221X1 U1331 (.IN1(n8), .IN2(n1281), .IN3(n1282), .IN4(n64), .IN5(n1283), .Q(n1247));
   AO22X1 U1332 (.IN1(n250), .IN2(n32), .IN3(n206), .IN4(n273), .Q(n1283));
   NAND4X0 U1333 (.IN1(n1266), .IN2(n53), .IN3(n203), .IN4(n1284), .QN(n1282));
   OA222X1 U1334 (.IN1(n225), .IN2(n38), .IN3(n7), .IN4(n56), .IN5(n49), .IN6(n1409), .Q(
          n1284));
   NAND3X0 U1335 (.IN1(n270), .IN2(n190), .IN3(n1286), .QN(n1281));
   AO222X1 U1336 (.IN1(n1210), .IN2(n1287), .IN3(n1212), .IN4(n1288), .IN5(sboxw[15]), .
          IN6(n1289), .Q(new_sboxw[12]));
   AO221X1 U1337 (.IN1(n177), .IN2(n1290), .IN3(n179), .IN4(n1291), .IN5(n1292), .Q(n1289)
          );
   AO22X1 U1338 (.IN1(n182), .IN2(n1293), .IN3(n184), .IN4(n1294), .Q(n1292));
   NAND4X0 U1339 (.IN1(n45), .IN2(n1232), .IN3(n1277), .IN4(n1295), .QN(n1294));
   OA222X1 U1340 (.IN1(n37), .IN2(n1413), .IN3(n194), .IN4(n1231), .IN5(n58), .IN6(n32), .
          Q(n1295));
   NAND4X0 U1341 (.IN1(n1297), .IN2(n190), .IN3(n1298), .IN4(n1299), .QN(n1293));
   OA222X1 U1342 (.IN1(n7), .IN2(n46), .IN3(n188), .IN4(n41), .IN5(n219), .IN6(n38), .Q(
          n1299));
   NAND4X0 U1343 (.IN1(n248), .IN2(n1266), .IN3(n1301), .IN4(n1302), .QN(n1291));
   OA222X1 U1344 (.IN1(n225), .IN2(n38), .IN3(n1303), .IN4(n1410), .IN5(n1415), .IN6(n37)
          , .Q(n1302));
   AO21X1 U1345 (.IN1(n43), .IN2(n53), .IN3(n1), .Q(n1301));
   OA221X1 U1346 (.IN1(n225), .IN2(n51), .IN3(n219), .IN4(n49), .IN5(n1261), .Q(n1305));
   OA222X1 U1347 (.IN1(n1415), .IN2(n213), .IN3(n6), .IN4(n41), .IN5(n7), .IN6(n47), .Q(
          n1304));
   AO222X1 U1348 (.IN1(n1306), .IN2(n64), .IN3(n8), .IN4(n1307), .IN5(n238), .IN6(n206), .
          Q(n1288));
   NAND4X0 U1349 (.IN1(n40), .IN2(n53), .IN3(n1205), .IN4(n1308), .QN(n1307));
   OA22X1 U1350 (.IN1(n1296), .IN2(n57), .IN3(n37), .IN4(n1411), .Q(n1308));
   NAND4X0 U1351 (.IN1(n210), .IN2(n1309), .IN3(n1310), .IN4(n1311), .QN(n1306));
   OA222X1 U1352 (.IN1(n6), .IN2(n60), .IN3(n194), .IN4(n38), .IN5(n1410), .IN6(n53), .Q(
          n1311));
   AO222X1 U1353 (.IN1(n206), .IN2(n39), .IN3(n8), .IN4(n1312), .IN5(n1313), .IN6(n64), .Q(
          n1287));
   NAND4X0 U1354 (.IN1(n40), .IN2(n1297), .IN3(n1314), .IN4(n1315), .QN(n1313));
   OA221X1 U1355 (.IN1(n1415), .IN2(n37), .IN3(n193), .IN4(n244), .IN5(n1316), .Q(n1315)
          );
   AND2X1 U1356 (.IN1(n1219), .IN2(n264), .Q(n1314));
   NAND4X0 U1357 (.IN1(n227), .IN2(n264), .IN3(n1300), .IN4(n1317), .QN(n1312));
   OA22X1 U1358 (.IN1(n1296), .IN2(n58), .IN3(n47), .IN4(n1409), .Q(n1317));
   OA22X1 U1359 (.IN1(n1409), .IN2(n48), .IN3(n1), .IN4(sboxw[10]), .Q(n1296));
   AO22X1 U1360 (.IN1(sboxw[15]), .IN2(n1319), .IN3(n1320), .IN4(n66), .Q(new_sboxw[11])
          );
   AO222X1 U1361 (.IN1(n179), .IN2(n1321), .IN3(n177), .IN4(n1322), .IN5(n1323), .IN6(n65)
          , .Q(n1320));
   AO222X1 U1362 (.IN1(n206), .IN2(n36), .IN3(n8), .IN4(n1324), .IN5(n1325), .IN6(n64), .Q(
          n1323));
   NAND4X0 U1363 (.IN1(n1300), .IN2(n1309), .IN3(n1326), .IN4(n1327), .QN(n1325));
   AND4X1 U1364 (.IN1(n1261), .IN2(n1266), .IN3(n1218), .IN4(n1182), .Q(n1327));
   NAND4X0 U1365 (.IN1(n1328), .IN2(n52), .IN3(n1203), .IN4(n1261), .QN(n1324));
   OR2X1 U1366 (.IN1(n1412), .IN2(n200), .Q(n1328));
   NAND4X0 U1367 (.IN1(n248), .IN2(n47), .IN3(n52), .IN4(n1329), .QN(n1322));
   OA222X1 U1368 (.IN1(n6), .IN2(n60), .IN3(n225), .IN4(n1330), .IN5(n200), .IN6(n1413), .
          Q(n1329));
   NAND4X0 U1369 (.IN1(n210), .IN2(n1331), .IN3(n1332), .IN4(n1333), .QN(n1321));
   AND4X1 U1370 (.IN1(n190), .IN2(n1266), .IN3(n216), .IN4(n1182), .Q(n1333));
   OA22X1 U1371 (.IN1(n1413), .IN2(n38), .IN3(n1414), .IN4(n46), .Q(n1332));
   AO222X1 U1372 (.IN1(n182), .IN2(n1334), .IN3(n184), .IN4(n1335), .IN5(sboxw[14]), .IN6(
          n1336), .Q(n1319));
   AO222X1 U1373 (.IN1(n261), .IN2(n206), .IN3(n8), .IN4(n1337), .IN5(n1338), .IN6(n64), .
          Q(n1336));
   NAND4X0 U1374 (.IN1(n1297), .IN2(n1218), .IN3(n1339), .IN4(n1340), .QN(n1338));
   OA222X1 U1375 (.IN1(n37), .IN2(n1413), .IN3(n1270), .IN4(n1415), .IN5(n57), .IN6(n1411)
          , .Q(n1340));
   AO21X1 U1376 (.IN1(n43), .IN2(n47), .IN3(n193), .Q(n1339));
   NAND4X0 U1377 (.IN1(n1331), .IN2(n1316), .IN3(n1341), .IN4(n1342), .QN(n1337));
   OA221X1 U1378 (.IN1(n213), .IN2(n1409), .IN3(n42), .IN4(n1414), .IN5(n214), .Q(n1342)
          );
   NAND4X0 U1379 (.IN1(n189), .IN2(n1219), .IN3(n1343), .IN4(n1344), .QN(n1335));
   OA222X1 U1380 (.IN1(n188), .IN2(n42), .IN3(n219), .IN4(n33), .IN5(n193), .IN6(n51), .Q(
          n1344));
   OR2X1 U1381 (.IN1(n1), .IN2(n1345), .Q(n1343));
   NAND4X0 U1382 (.IN1(n270), .IN2(n248), .IN3(n1346), .IN4(n1347), .QN(n1334));
   OA22X1 U1383 (.IN1(n1413), .IN2(n53), .IN3(n1412), .IN4(n43), .Q(n1347));
   AO222X1 U1384 (.IN1(n172), .IN2(n1348), .IN3(n174), .IN4(n1349), .IN5(n1350), .IN6(n66)
          , .Q(new_sboxw[10]));
   AO222X1 U1385 (.IN1(n182), .IN2(n1351), .IN3(n184), .IN4(n1352), .IN5(sboxw[14]), .IN6(
          n1353), .Q(n1350));
   NAND4X0 U1386 (.IN1(n1203), .IN2(n190), .IN3(n1354), .IN4(n1355), .QN(n1353));
   OA22X1 U1387 (.IN1(n8), .IN2(n1356), .IN3(n63), .IN4(n37), .Q(n1355));
   NOR4X0 U1388 (.IN1(n1357), .IN2(n1358), .IN3(n269), .IN4(n1245), .QN(n1356));
   AO222X1 U1389 (.IN1(n225), .IN2(n261), .IN3(n240), .IN4(n1415), .IN5(sboxw[11]), .IN6(
          n1411), .Q(n1357));
   NAND3X0 U1390 (.IN1(n1232), .IN2(n216), .IN3(n202), .QN(n1359));
   NAND4X0 U1391 (.IN1(n1316), .IN2(n196), .IN3(n1360), .IN4(n1361), .QN(n1352));
   AND2X1 U1392 (.IN1(n255), .IN2(n1179), .Q(n1361));
   OA22X1 U1393 (.IN1(n47), .IN2(n1414), .IN3(n38), .IN4(n1411), .Q(n255));
   NAND4X0 U1394 (.IN1(n1309), .IN2(n227), .IN3(n1362), .IN4(n1363), .QN(n1351));
   OA221X1 U1395 (.IN1(n1411), .IN2(n53), .IN3(n194), .IN4(n47), .IN5(n1187), .Q(n1363));
   OA22X1 U1396 (.IN1(n7), .IN2(n41), .IN3(n1414), .IN4(n38), .Q(n1362));
   AO22X1 U1397 (.IN1(n8), .IN2(n1364), .IN3(n1365), .IN4(n64), .Q(n1349));
   NAND4X0 U1398 (.IN1(n1183), .IN2(n35), .IN3(n1366), .IN4(n1367), .QN(n1365));
   OA22X1 U1399 (.IN1(n1414), .IN2(n58), .IN3(n193), .IN4(n46), .Q(n1367));
   NAND4X0 U1400 (.IN1(n1277), .IN2(n1181), .IN3(n1368), .IN4(n1369), .QN(n1364));
   OA222X1 U1401 (.IN1(n1414), .IN2(n38), .IN3(n1345), .IN4(n1413), .IN5(n41), .IN6(n1412)
          , .Q(n1369));
   AND2X1 U1402 (.IN1(n1203), .IN2(n224), .Q(n1368));
   AO22X1 U1403 (.IN1(n8), .IN2(n1370), .IN3(n1371), .IN4(n64), .Q(n1348));
   NAND4X0 U1404 (.IN1(n1205), .IN2(n1331), .IN3(n1372), .IN4(n1373), .QN(n1371));
   OA222X1 U1405 (.IN1(n7), .IN2(n53), .IN3(n51), .IN4(n1414), .IN5(n193), .IN6(n38), .Q(
          n1373));
   AND2X1 U1406 (.IN1(n1219), .IN2(n227), .Q(n1372));
   AO221X1 U1407 (.IN1(n205), .IN2(n1413), .IN3(n238), .IN4(n219), .IN5(n1374), .Q(n1370)
          );
   OAI221X1 U1408 (.IN1(n1411), .IN2(n49), .IN3(n1303), .IN4(n193), .IN5(n1181), .QN(n1374)
          );
   AO222X1 U1409 (.IN1(n598), .IN2(n1375), .IN3(n600), .IN4(n1376), .IN5(n1377), .IN6(
          n1408), .Q(new_sboxw[0]));
   AO222X1 U1410 (.IN1(n308), .IN2(n1378), .IN3(n310), .IN4(n1379), .IN5(sboxw[6]), .IN6(
          n1380), .Q(n1377));
   AO221X1 U1411 (.IN1(n1381), .IN2(n14), .IN3(n13), .IN4(n1382), .IN5(n495), .Q(n1380));
   NAND4X0 U1412 (.IN1(n286), .IN2(n153), .IN3(n1383), .IN4(n1384), .QN(n1382));
   OA222X1 U1413 (.IN1(n401), .IN2(n26), .IN3(n302), .IN4(n171), .IN5(n1404), .IN6(n29), .
          Q(n1384));
   AO22X1 U1414 (.IN1(n335), .IN2(n106), .IN3(n476), .IN4(n22), .Q(n1381));
   NAND4X0 U1415 (.IN1(n290), .IN2(n1385), .IN3(n1386), .IN4(n440), .QN(n1379));
   OR2X1 U1416 (.IN1(n1404), .IN2(n297), .Q(n1385));
   OA22X1 U1417 (.IN1(n163), .IN2(n106), .IN3(n25), .IN4(sboxw[2]), .Q(n297));
   OA221X1 U1418 (.IN1(n160), .IN2(n25), .IN3(n171), .IN4(n27), .IN5(n157), .Q(n290));
   NAND4X0 U1419 (.IN1(n322), .IN2(n362), .IN3(n1387), .IN4(n1388), .QN(n1378));
   OA221X1 U1420 (.IN1(n288), .IN2(n1405), .IN3(n4), .IN4(n1402), .IN5(n456), .Q(n1388));
   OR2X1 U1421 (.IN1(n29), .IN2(n394), .Q(n1387));
   NAND3X0 U1422 (.IN1(n615), .IN2(n1389), .IN3(n1390), .QN(n1376));
   OA222X1 U1423 (.IN1(n152), .IN2(n107), .IN3(n13), .IN4(n1391), .IN5(n1392), .IN6(n14), .
          Q(n1390));
   OA221X1 U1424 (.IN1(n302), .IN2(n1404), .IN3(n25), .IN4(n171), .IN5(n1393), .Q(n1392)
          );
   OA221X1 U1425 (.IN1(n319), .IN2(n164), .IN3(n288), .IN4(n171), .IN5(n1394), .Q(n1391)
          );
   AND2X1 U1426 (.IN1(n154), .IN2(n325), .Q(n1394));
   OA22X1 U1427 (.IN1(n154), .IN2(n29), .IN3(n158), .IN4(n22), .Q(n615));
   AO221X1 U1428 (.IN1(n1395), .IN2(n14), .IN3(n13), .IN4(n1396), .IN5(n1397), .Q(n1375)
          );
   AO22X1 U1429 (.IN1(n470), .IN2(n281), .IN3(n305), .IN4(n29), .Q(n1397));
   NAND4X0 U1430 (.IN1(n424), .IN2(n158), .IN3(n1398), .IN4(n1399), .QN(n1396));
   OA22X1 U1431 (.IN1(n288), .IN2(n1402), .IN3(n106), .IN4(n164), .Q(n1399));
   AO221X1 U1432 (.IN1(n288), .IN2(n303), .IN3(n291), .IN4(n30), .IN5(n1400), .Q(n1395));
   AO21X1 U1433 (.IN1(n1401), .IN2(n29), .IN3(n1043), .Q(n1400));
   NBUFFX2 U1 (.INP(sboxw[24]), .Z(n11));
   NBUFFX2 U2 (.INP(sboxw[16]), .Z(n9));
   NBUFFX2 U3 (.INP(sboxw[0]), .Z(n4));
   NBUFFX2 U4 (.INP(sboxw[8]), .Z(n6));
   NBUFFX2 U5 (.INP(sboxw[9]), .Z(n7));
   NBUFFX2 U6 (.INP(sboxw[13]), .Z(n8));
   INVX0 U7 (.INP(n316), .ZN(n28));
   INVX0 U8 (.INP(n878), .ZN(n77));
   INVX0 U9 (.INP(n1112), .ZN(n69));
   INVX0 U10 (.INP(n625), .ZN(n20));
   INVX0 U11 (.INP(n777), .ZN(n113));
   NOR2X0 U12 (.IN1(n29), .IN2(n157), .QN(n316));
   NOR2X0 U13 (.IN1(n78), .IN2(n89), .QN(n878));
   NAND2X1 U14 (.IN1(n131), .IN2(n119), .QN(n819));
   NOR2X0 U15 (.IN1(n71), .IN2(n85), .QN(n1112));
   NOR2X0 U16 (.IN1(n22), .IN2(n153), .QN(n625));
   NOR2X0 U17 (.IN1(n115), .IN2(n129), .QN(n777));
   INVX0 U18 (.INP(n1242), .ZN(n52));
   INVX0 U19 (.INP(n536), .ZN(n121));
   INVX0 U20 (.INP(n1190), .ZN(n45));
   INVX0 U21 (.INP(n1200), .ZN(n40));
   NAND2X1 U22 (.IN1(n37), .IN2(n41), .QN(n1258));
   NAND2X1 U23 (.IN1(n869), .IN2(n78), .QN(n907));
   NAND2X1 U24 (.IN1(n307), .IN2(n29), .QN(n345));
   OA21X1 U25 (.IN1(n165), .IN2(n30), .IN3(n345), .Q(n298));
   OA21X1 U26 (.IN1(n97), .IN2(n79), .IN3(n907), .Q(n860));
   NAND2X1 U27 (.IN1(n291), .IN2(n29), .QN(n449));
   NAND2X1 U28 (.IN1(n853), .IN2(n78), .QN(n1011));
   OA21X1 U29 (.IN1(n29), .IN2(n151), .IN3(n439), .Q(n437));
   OA21X1 U30 (.IN1(n78), .IN2(n83), .IN3(n1001), .Q(n999));
   NAND3X0 U31 (.IN1(n554), .IN2(n3), .IN3(n674), .QN(n592));
   INVX0 U32 (.INP(n288), .ZN(n26));
   NAND2X1 U33 (.IN1(n307), .IN2(n26), .QN(n356));
   INVX0 U34 (.INP(n850), .ZN(n75));
   NAND2X1 U35 (.IN1(n869), .IN2(n75), .QN(n918));
   NAND2X1 U36 (.IN1(n1069), .IN2(n75), .QN(n925));
   INVX0 U37 (.INP(n508), .ZN(n119));
   NAND2X1 U38 (.IN1(n527), .IN2(n119), .QN(n576));
   NAND2X1 U39 (.IN1(n480), .IN2(n26), .QN(n363));
   NAND2X1 U40 (.IN1(n734), .IN2(n119), .QN(n583));
   NAND2X1 U41 (.IN1(n291), .IN2(n26), .QN(n458));
   NAND2X1 U42 (.IN1(n853), .IN2(n75), .QN(n1020));
   NAND2X1 U43 (.IN1(n511), .IN2(n119), .QN(n712));
   INVX0 U44 (.INP(n225), .ZN(n1410));
   NAND2X1 U45 (.IN1(n239), .IN2(n1410), .QN(n1183));
   INVX0 U46 (.INP(n896), .ZN(n71));
   NOR2X0 U47 (.IN1(n97), .IN2(n71), .QN(n882));
   NOR2X0 U48 (.IN1(n853), .IN2(n882), .QN(n1164));
   NAND2X1 U49 (.IN1(n238), .IN2(n1410), .QN(n190));
   INVX0 U50 (.INP(n334), .ZN(n22));
   NOR2X0 U51 (.IN1(n165), .IN2(n22), .QN(n320));
   NOR2X0 U52 (.IN1(n291), .IN2(n320), .QN(n1393));
   NAND2X1 U53 (.IN1(n205), .IN2(n1410), .QN(n1232));
   NAND2X1 U54 (.IN1(n480), .IN2(n22), .QN(n400));
   OA21X1 U55 (.IN1(n25), .IN2(n167), .IN3(n423), .Q(n422));
   OA21X1 U56 (.IN1(n158), .IN2(n288), .IN3(n400), .Q(n423));
   NAND2X1 U57 (.IN1(n1069), .IN2(n71), .QN(n962));
   OA21X1 U58 (.IN1(n74), .IN2(n99), .IN3(n985), .Q(n984));
   OA21X1 U59 (.IN1(n90), .IN2(n850), .IN3(n962), .Q(n985));
   INVX0 U60 (.INP(n554), .ZN(n115));
   NOR2X0 U61 (.IN1(n141), .IN2(n115), .QN(n540));
   NOR2X0 U62 (.IN1(n511), .IN2(n540), .QN(n829));
   NAND2X1 U63 (.IN1(n734), .IN2(n115), .QN(n654));
   OA21X1 U64 (.IN1(n134), .IN2(n508), .IN3(n654), .Q(n677));
   OA21X1 U65 (.IN1(n118), .IN2(n143), .IN3(n677), .Q(n676));
   NAND2X1 U66 (.IN1(n261), .IN2(n1410), .QN(n227));
   NAND2X1 U67 (.IN1(n288), .IN2(n420), .QN(n405));
   NAND2X1 U68 (.IN1(n850), .IN2(n982), .QN(n967));
   NAND2X1 U69 (.IN1(n188), .IN2(n1285), .QN(n1286));
   OA21X1 U70 (.IN1(n164), .IN2(n288), .IN3(n400), .Q(n468));
   OA21X1 U71 (.IN1(n96), .IN2(n850), .IN3(n962), .Q(n1057));
   NAND2X1 U72 (.IN1(n508), .IN2(n674), .QN(n659));
   OA21X1 U73 (.IN1(n140), .IN2(n508), .IN3(n654), .Q(n722));
   NOR2X0 U74 (.IN1(n1409), .IN2(n53), .QN(n1242));
   NOR2X0 U75 (.IN1(n2), .IN2(n133), .QN(n536));
   INVX0 U76 (.INP(n188), .ZN(n1411));
   NOR2X0 U77 (.IN1(n1411), .IN2(n51), .QN(n262));
   NOR2X0 U78 (.IN1(n261), .IN2(n262), .QN(n260));
   OA21X1 U79 (.IN1(n850), .IN2(n851), .IN3(n852), .Q(n849));
   NAND2X1 U80 (.IN1(n527), .IN2(n2), .QN(n565));
   NOR2X0 U81 (.IN1(n1409), .IN2(n46), .QN(n1190));
   OA21X1 U82 (.IN1(n141), .IN2(n123), .IN3(n565), .Q(n518));
   NAND2X1 U83 (.IN1(n205), .IN2(n1411), .QN(n1266));
   NOR2X0 U84 (.IN1(n41), .IN2(n1), .QN(n1200));
   NAND2X1 U85 (.IN1(n238), .IN2(n1), .QN(n1219));
   OA21X1 U86 (.IN1(n1413), .IN2(n51), .IN3(n1219), .Q(n1187));
   NAND2X1 U87 (.IN1(n1258), .IN2(n1409), .QN(n1346));
   NAND2X1 U88 (.IN1(n511), .IN2(n2), .QN(n703));
   NAND2X1 U89 (.IN1(n420), .IN2(n30), .QN(n344));
   NAND2X1 U90 (.IN1(n982), .IN2(n79), .QN(n906));
   NAND2X1 U91 (.IN1(n674), .IN2(n123), .QN(n564));
   INVX0 U92 (.INP(n1140), .ZN(n80));
   INVX0 U93 (.INP(n1043), .ZN(n31));
   OA21X1 U94 (.IN1(n122), .IN2(n127), .IN3(n693), .Q(n691));
   NAND2X1 U95 (.IN1(n896), .IN2(n926), .QN(n920));
   NAND2X1 U96 (.IN1(n334), .IN2(n364), .QN(n358));
   OA21X1 U97 (.IN1(n154), .IN2(n30), .IN3(n152), .Q(n490));
   OA21X1 U98 (.IN1(n86), .IN2(n79), .IN3(n84), .Q(n1079));
   NAND2X1 U99 (.IN1(n554), .IN2(n584), .QN(n578));
   INVX0 U100 (.INP(n805), .ZN(n124));
   OA21X1 U101 (.IN1(n130), .IN2(n123), .IN3(n128), .Q(n744));
   NOR2X0 U102 (.IN1(n55), .IN2(n1413), .QN(n1245));
   NAND2X1 U103 (.IN1(n1285), .IN2(n1413), .QN(n1218));
   NAND2X1 U104 (.IN1(n261), .IN2(n1), .QN(n210));
   OA21X1 U105 (.IN1(n1414), .IN2(n34), .IN3(n1300), .Q(n1298));
   NAND2X1 U106 (.IN1(n238), .IN2(n188), .QN(n224));
   NAND2X1 U107 (.IN1(n188), .IN2(n1258), .QN(n1255));
   INVX0 U108 (.INP(n495), .ZN(n18));
   INVX0 U109 (.INP(n1084), .ZN(n67));
   OA21X1 U110 (.IN1(n1413), .IN2(n47), .IN3(n46), .Q(n214));
   INVX0 U111 (.INP(n749), .ZN(n111));
   OA21X1 U112 (.IN1(n46), .IN2(n188), .IN3(n1274), .Q(n1179));
   NAND2X1 U113 (.IN1(n140), .IN2(n134), .QN(n689));
   NAND2X1 U114 (.IN1(n96), .IN2(n90), .QN(n997));
   NAND2X1 U115 (.IN1(n91), .IN2(n97), .QN(n926));
   INVX0 U116 (.INP(n261), .ZN(n37));
   NAND2X1 U117 (.IN1(n135), .IN2(n141), .QN(n584));
   INVX0 U118 (.INP(n205), .ZN(n47));
   NAND2X1 U119 (.IN1(n164), .IN2(n158), .QN(n435));
   INVX0 U120 (.INP(n1069), .ZN(n86));
   INVX0 U121 (.INP(n734), .ZN(n130));
   INVX0 U122 (.INP(n1018), .ZN(n87));
   NAND2X1 U123 (.IN1(n159), .IN2(n165), .QN(n364));
   INVX0 U124 (.INP(n710), .ZN(n131));
   INVX0 U125 (.INP(n1285), .ZN(n41));
   INVX0 U126 (.INP(n239), .ZN(n42));
   INVX0 U127 (.INP(n511), .ZN(n138));
   INVX0 U128 (.INP(n853), .ZN(n94));
   NOR2X0 U129 (.IN1(n511), .IN2(n674), .QN(n645));
   NOR2X0 U130 (.IN1(n853), .IN2(n982), .QN(n953));
   INVX0 U131 (.INP(n555), .ZN(n135));
   INVX0 U132 (.INP(n674), .ZN(n133));
   INVX0 U133 (.INP(n335), .ZN(n159));
   INVX0 U134 (.INP(n420), .ZN(n157));
   INVX0 U135 (.INP(n480), .ZN(n154));
   INVX0 U136 (.INP(n897), .ZN(n91));
   INVX0 U137 (.INP(n982), .ZN(n89));
   INVX0 U138 (.INP(n869), .ZN(n85));
   INVX0 U139 (.INP(n238), .ZN(n43));
   NAND2X1 U140 (.IN1(n61), .IN2(n43), .QN(n1201));
   INVX0 U141 (.INP(n527), .ZN(n129));
   INVX0 U142 (.INP(n456), .ZN(n155));
   INVX0 U143 (.INP(n291), .ZN(n162));
   NOR2X0 U144 (.IN1(n291), .IN2(n420), .QN(n391));
   INVX0 U145 (.INP(n1231), .ZN(n39));
   INVX0 U146 (.INP(n307), .ZN(n153));
   NAND2X1 U147 (.IN1(n1404), .IN2(n153), .QN(n317));
   NAND2X1 U148 (.IN1(n105), .IN2(n83), .QN(n1109));
   NAND2X1 U149 (.IN1(n60), .IN2(n34), .QN(n201));
   NAND2X1 U150 (.IN1(n149), .IN2(n127), .QN(n774));
   NAND2X1 U151 (.IN1(n1405), .IN2(n151), .QN(n622));
   INVX0 U152 (.INP(n1065), .ZN(n92));
   INVX0 U153 (.INP(n240), .ZN(n35));
   INVX0 U154 (.INP(n730), .ZN(n136));
   INVX0 U155 (.INP(n476), .ZN(n160));
   INVX0 U156 (.INP(n269), .ZN(n58));
   INVX0 U157 (.INP(n525), .ZN(n145));
   INVX0 U158 (.INP(n867), .ZN(n101));
   INVX0 U159 (.INP(n305), .ZN(n171));
   NOR2X0 U160 (.IN1(n109), .IN2(n15), .QN(n948));
   NAND2X1 U161 (.IN1(n15), .IN2(n1098), .QN(n1093));
   NOR2X0 U162 (.IN1(n1096), .IN2(n1097), .QN(n1095));
   NAND2X1 U163 (.IN1(n975), .IN2(n864), .QN(n970));
   NAND2X1 U164 (.IN1(n413), .IN2(n302), .QN(n408));
   NAND2X1 U165 (.IN1(n413), .IN2(n27), .QN(n1041));
   NAND2X1 U166 (.IN1(n975), .IN2(n76), .QN(n1138));
   NAND2X1 U167 (.IN1(n1105), .IN2(n78), .QN(n883));
   NAND2X1 U168 (.IN1(n618), .IN2(n29), .QN(n321));
   NOR2X0 U169 (.IN1(n854), .IN2(n68), .QN(n1101));
   INVX0 U170 (.INP(n1102), .ZN(n68));
   NOR2X0 U171 (.IN1(n292), .IN2(n19), .QN(n614));
   INVX0 U172 (.INP(n615), .ZN(n19));
   NAND2X1 U173 (.IN1(n333), .IN2(n29), .QN(n365));
   NAND2X1 U174 (.IN1(n895), .IN2(n78), .QN(n927));
   NAND2X1 U175 (.IN1(n13), .IN2(n611), .QN(n606));
   NOR2X0 U176 (.IN1(n609), .IN2(n610), .QN(n608));
   INVX0 U177 (.INP(n425), .ZN(n24));
   INVX0 U178 (.INP(n987), .ZN(n73));
   NAND2X1 U179 (.IN1(n975), .IN2(n896), .QN(n1117));
   NAND2X1 U180 (.IN1(n164), .IN2(n160), .QN(n1401));
   NAND2X1 U181 (.IN1(n413), .IN2(n334), .QN(n630));
   NAND2X1 U182 (.IN1(n96), .IN2(n92), .QN(n1172));
   INVX0 U183 (.INP(n17), .ZN(n3));
   INVX0 U184 (.INP(n843), .ZN(n82));
   NOR2X0 U185 (.IN1(n1407), .IN2(n13), .QN(n386));
   NOR2X0 U186 (.IN1(n302), .IN2(n328), .QN(n288));
   NOR2X0 U187 (.IN1(n864), .IN2(n890), .QN(n850));
   NOR2X0 U188 (.IN1(n522), .IN2(n548), .QN(n508));
   NOR2X0 U189 (.IN1(n193), .IN2(n219), .QN(n225));
   NOR2X0 U190 (.IN1(n81), .IN2(n76), .QN(n896));
   NOR2X0 U191 (.IN1(n106), .IN2(n27), .QN(n334));
   NAND2X1 U192 (.IN1(n1318), .IN2(n1410), .QN(n1182));
   NOR2X0 U193 (.IN1(n125), .IN2(n120), .QN(n554));
   NAND2X1 U194 (.IN1(n288), .IN2(n303), .QN(n491));
   INVX0 U195 (.INP(n333), .ZN(n168));
   NAND2X1 U196 (.IN1(n850), .IN2(n865), .QN(n1080));
   INVX0 U197 (.INP(n895), .ZN(n100));
   NAND2X1 U198 (.IN1(n104), .IN2(n85), .QN(n879));
   NAND2X1 U199 (.IN1(n508), .IN2(n523), .QN(n745));
   INVX0 U200 (.INP(n553), .ZN(n144));
   NAND2X1 U201 (.IN1(n288), .IN2(n618), .QN(n448));
   NAND2X1 U202 (.IN1(n850), .IN2(n1105), .QN(n1010));
   NAND2X1 U203 (.IN1(n148), .IN2(n129), .QN(n537));
   NAND2X1 U204 (.IN1(n508), .IN2(n770), .QN(n702));
   NOR2X0 U205 (.IN1(n512), .IN2(n112), .QN(n766));
   INVX0 U206 (.INP(n767), .ZN(n112));
   NAND2X1 U207 (.IN1(n201), .IN2(n1411), .QN(n1366));
   INVX0 U208 (.INP(n193), .ZN(n1409));
   NAND2X1 U209 (.IN1(n1059), .IN2(n71), .QN(n974));
   INVX0 U210 (.INP(n328), .ZN(n25));
   NAND2X1 U211 (.IN1(n470), .IN2(n25), .QN(n388));
   INVX0 U212 (.INP(n890), .ZN(n74));
   NAND2X1 U213 (.IN1(n1059), .IN2(n74), .QN(n950));
   NAND2X1 U214 (.IN1(n225), .IN2(n273), .QN(n189));
   NAND2X1 U215 (.IN1(n470), .IN2(n22), .QN(n412));
   INVX0 U216 (.INP(n548), .ZN(n118));
   NAND2X1 U217 (.IN1(n724), .IN2(n118), .QN(n642));
   NOR2X0 U218 (.IN1(n1412), .IN2(n1415), .QN(n188));
   NOR2X0 U219 (.IN1(n330), .IN2(n335), .QN(n399));
   NOR2X0 U220 (.IN1(n892), .IN2(n897), .QN(n961));
   NAND2X1 U221 (.IN1(n280), .IN2(n22), .QN(n436));
   NAND2X1 U222 (.IN1(n842), .IN2(n71), .QN(n998));
   NAND2X1 U223 (.IN1(n724), .IN2(n115), .QN(n666));
   NAND2X1 U224 (.IN1(n667), .IN2(n522), .QN(n662));
   NOR2X0 U225 (.IN1(n550), .IN2(n555), .QN(n653));
   NAND2X1 U226 (.IN1(n500), .IN2(n115), .QN(n690));
   NAND2X1 U227 (.IN1(n667), .IN2(n554), .QN(n782));
   NAND2X1 U228 (.IN1(n330), .IN2(n302), .QN(n1398));
   NAND2X1 U229 (.IN1(n892), .IN2(n864), .QN(n1169));
   NAND2X1 U230 (.IN1(n550), .IN2(n522), .QN(n834));
   NAND2X1 U231 (.IN1(n1280), .IN2(n225), .QN(n1309));
   INVX0 U232 (.INP(n1296), .ZN(n32));
   NAND2X1 U233 (.IN1(n302), .IN2(n364), .QN(n1386));
   NAND2X1 U234 (.IN1(n864), .IN2(n926), .QN(n1157));
   NAND2X1 U235 (.IN1(n140), .IN2(n136), .QN(n837));
   NAND2X1 U236 (.IN1(n667), .IN2(n120), .QN(n803));
   NAND2X1 U237 (.IN1(n522), .IN2(n584), .QN(n822));
   NAND2X1 U238 (.IN1(n770), .IN2(n122), .QN(n541));
   NAND2X1 U239 (.IN1(n328), .IN2(n318), .QN(n424));
   NAND2X1 U240 (.IN1(n890), .IN2(n880), .QN(n986));
   NAND2X1 U241 (.IN1(n268), .IN2(n1411), .QN(n1277));
   NAND2X1 U242 (.IN1(n215), .IN2(n219), .QN(n1273));
   NAND2X1 U243 (.IN1(n225), .IN2(n1258), .QN(n1360));
   NOR2X0 U244 (.IN1(n221), .IN2(n239), .QN(n1265));
   NAND2X1 U245 (.IN1(n160), .IN2(n1402), .QN(n332));
   NAND2X1 U246 (.IN1(n1318), .IN2(n1411), .QN(n1297));
   NAND2X1 U247 (.IN1(n92), .IN2(n102), .QN(n894));
   NAND2X1 U248 (.IN1(n136), .IN2(n146), .QN(n552));
   INVX0 U249 (.INP(n679), .ZN(n117));
   NAND2X1 U250 (.IN1(n864), .IN2(n853), .QN(n919));
   NAND2X1 U251 (.IN1(n548), .IN2(n538), .QN(n678));
   NAND2X1 U252 (.IN1(n330), .IN2(n334), .QN(n395));
   NAND2X1 U253 (.IN1(n892), .IN2(n896), .QN(n957));
   NAND2X1 U254 (.IN1(n302), .IN2(n291), .QN(n357));
   NAND2X1 U255 (.IN1(n522), .IN2(n511), .QN(n577));
   OA21X1 U256 (.IN1(n1414), .IN2(n53), .IN3(n47), .Q(n226));
   NAND2X1 U257 (.IN1(n328), .IN2(n618), .QN(n294));
   NAND2X1 U258 (.IN1(n550), .IN2(n554), .QN(n649));
   NAND2X1 U259 (.IN1(n890), .IN2(n1105), .QN(n856));
   INVX0 U260 (.INP(n319), .ZN(n30));
   INVX0 U261 (.INP(n881), .ZN(n79));
   NAND2X1 U262 (.IN1(n221), .IN2(n219), .QN(n271));
   NAND2X1 U263 (.IN1(n548), .IN2(n770), .QN(n514));
   INVX0 U264 (.INP(n539), .ZN(n123));
   NAND2X1 U265 (.IN1(n890), .IN2(n842), .QN(n913));
   NOR2X0 U266 (.IN1(n97), .IN2(n881), .QN(n1140));
   NOR2X0 U267 (.IN1(n165), .IN2(n319), .QN(n1043));
   NAND2X1 U268 (.IN1(n328), .IN2(n280), .QN(n351));
   NAND2X1 U269 (.IN1(n553), .IN2(n2), .QN(n585));
   NAND2X1 U270 (.IN1(n275), .IN2(n216), .QN(n274));
   NAND2X1 U271 (.IN1(n329), .IN2(n334), .QN(n286));
   NAND2X1 U272 (.IN1(n891), .IN2(n896), .QN(n848));
   NAND2X1 U273 (.IN1(n548), .IN2(n500), .QN(n571));
   NAND2X1 U274 (.IN1(n328), .IN2(n307), .QN(n467));
   NAND2X1 U275 (.IN1(n890), .IN2(n869), .QN(n1056));
   NAND2X1 U276 (.IN1(n549), .IN2(n554), .QN(n506));
   NAND2X1 U277 (.IN1(n548), .IN2(n527), .QN(n721));
   NAND2X1 U278 (.IN1(n35), .IN2(n57), .QN(n1209));
   NAND2X1 U279 (.IN1(n215), .IN2(n1412), .QN(n217));
   NOR2X0 U280 (.IN1(n141), .IN2(n539), .QN(n805));
   NAND2X1 U281 (.IN1(n250), .IN2(n251), .QN(n246));
   NAND2X1 U282 (.IN1(n1280), .IN2(n1414), .QN(n1203));
   NAND2X1 U283 (.IN1(n307), .IN2(n319), .QN(n409));
   NAND2X1 U284 (.IN1(n869), .IN2(n881), .QN(n971));
   INVX0 U285 (.INP(n1245), .ZN(n54));
   INVX0 U286 (.INP(n194), .ZN(n1413));
   NAND2X1 U287 (.IN1(n268), .IN2(n1413), .QN(n216));
   NAND2X1 U288 (.IN1(n1184), .IN2(n188), .QN(n241));
   NAND2X1 U289 (.IN1(n527), .IN2(n539), .QN(n663));
   NAND2X1 U290 (.IN1(n221), .IN2(n188), .QN(n1261));
   INVX0 U291 (.INP(n206), .ZN(n63));
   NAND2X1 U292 (.IN1(n193), .IN2(n238), .QN(n1326));
   NAND2X1 U293 (.IN1(n420), .IN2(n319), .QN(n359));
   NAND2X1 U294 (.IN1(n982), .IN2(n881), .QN(n921));
   NAND2X1 U295 (.IN1(n881), .IN2(n1105), .QN(n847));
   NAND2X1 U296 (.IN1(n319), .IN2(n618), .QN(n285));
   NAND2X1 U297 (.IN1(n193), .IN2(n1202), .QN(n270));
   NAND2X1 U298 (.IN1(n674), .IN2(n539), .QN(n579));
   NAND2X1 U299 (.IN1(n539), .IN2(n770), .QN(n505));
   NAND2X1 U300 (.IN1(n1207), .IN2(n1), .QN(n1233));
   NOR2X0 U301 (.IN1(n153), .IN2(n27), .QN(n495));
   NOR2X0 U302 (.IN1(n85), .IN2(n76), .QN(n1084));
   NOR2X0 U303 (.IN1(n129), .IN2(n120), .QN(n749));
   NAND2X1 U304 (.IN1(n1105), .IN2(n76), .QN(n887));
   NAND2X1 U305 (.IN1(n261), .IN2(n219), .QN(n1225));
   NAND2X1 U306 (.IN1(n618), .IN2(n27), .QN(n325));
   NOR2X0 U307 (.IN1(n65), .IN2(n64), .QN(n179));
   NAND2X1 U308 (.IN1(n280), .IN2(n27), .QN(n612));
   OA21X1 U309 (.IN1(n472), .IN2(n27), .IN3(n612), .Q(n1032));
   NAND2X1 U310 (.IN1(n842), .IN2(n76), .QN(n1099));
   OA21X1 U311 (.IN1(n1061), .IN2(n76), .IN3(n1099), .Q(n1129));
   NAND2X1 U312 (.IN1(n470), .IN2(n27), .QN(n439));
   NAND2X1 U313 (.IN1(n1059), .IN2(n76), .QN(n1001));
   NAND2X1 U314 (.IN1(n770), .IN2(n120), .QN(n545));
   OA21X1 U315 (.IN1(n152), .IN2(n319), .IN3(n162), .Q(n348));
   OA21X1 U316 (.IN1(n84), .IN2(n881), .IN3(n94), .Q(n910));
   NAND2X1 U317 (.IN1(n500), .IN2(n120), .QN(n764));
   OA21X1 U318 (.IN1(n726), .IN2(n120), .IN3(n764), .Q(n794));
   NAND2X1 U319 (.IN1(n724), .IN2(n120), .QN(n693));
   OA21X1 U320 (.IN1(n128), .IN2(n539), .IN3(n138), .Q(n568));
   NAND2X1 U321 (.IN1(n238), .IN2(n194), .QN(n1274));
   NAND2X1 U322 (.IN1(n333), .IN2(n106), .QN(n421));
   NAND2X1 U323 (.IN1(n895), .IN2(n81), .QN(n983));
   NAND2X1 U324 (.IN1(n291), .IN2(n27), .QN(n284));
   NAND2X1 U325 (.IN1(n853), .IN2(n76), .QN(n846));
   NAND2X1 U326 (.IN1(n1280), .IN2(n194), .QN(n197));
   NAND2X1 U327 (.IN1(n553), .IN2(n125), .QN(n675));
   NAND2X1 U328 (.IN1(n511), .IN2(n120), .QN(n504));
   NAND2X1 U329 (.IN1(n1280), .IN2(n1412), .QN(n264));
   NAND2X1 U330 (.IN1(n194), .IN2(n1285), .QN(n203));
   NAND2X1 U331 (.IN1(n1318), .IN2(n1412), .QN(n196));
   OA21X1 U332 (.IN1(n195), .IN2(n1412), .IN3(n196), .Q(n191));
   NAND2X1 U333 (.IN1(n268), .IN2(n1412), .QN(n1300));
   INVX0 U334 (.INP(n1318), .ZN(n53));
   INVX0 U335 (.INP(n250), .ZN(n61));
   NAND2X1 U336 (.IN1(n261), .IN2(n1412), .QN(n1181));
   NOR2X0 U337 (.IN1(n1415), .IN2(n49), .QN(n1358));
   INVX0 U338 (.INP(n1202), .ZN(n60));
   INVX0 U339 (.INP(n268), .ZN(n51));
   INVX0 U340 (.INP(n1059), .ZN(n97));
   INVX0 U341 (.INP(n880), .ZN(n105));
   INVX0 U342 (.INP(n281), .ZN(n107));
   OA21X1 U343 (.IN1(n46), .IN2(n194), .IN3(n37), .Q(n1222));
   NAND2X1 U344 (.IN1(n291), .IN2(n106), .QN(n1389));
   NAND2X1 U345 (.IN1(n853), .IN2(n81), .QN(n1160));
   INVX0 U346 (.INP(n501), .ZN(n126));
   INVX0 U347 (.INP(n500), .ZN(n140));
   INVX0 U348 (.INP(n670), .ZN(n148));
   INVX0 U349 (.INP(n842), .ZN(n96));
   INVX0 U350 (.INP(n978), .ZN(n104));
   INVX0 U351 (.INP(n724), .ZN(n141));
   INVX0 U352 (.INP(n538), .ZN(n149));
   NAND2X1 U353 (.IN1(n511), .IN2(n125), .QN(n825));
   NOR2X0 U354 (.IN1(n61), .IN2(n48), .QN(n261));
   NOR2X0 U355 (.IN1(n48), .IN2(n60), .QN(n205));
   INVX0 U356 (.INP(n280), .ZN(n164));
   NOR2X0 U357 (.IN1(n105), .IN2(n95), .QN(n1069));
   INVX0 U358 (.INP(n470), .ZN(n165));
   NOR2X0 U359 (.IN1(n149), .IN2(n139), .QN(n734));
   NOR2X0 U360 (.IN1(n1069), .IN2(n868), .QN(n1018));
   NOR2X0 U361 (.IN1(n734), .IN2(n526), .QN(n710));
   NOR2X0 U362 (.IN1(n239), .IN2(n268), .QN(n249));
   INVX0 U363 (.INP(n318), .ZN(n1405));
   NAND2X1 U364 (.IN1(n261), .IN2(n1415), .QN(n256));
   NOR2X0 U365 (.IN1(n1193), .IN2(n268), .QN(n1270));
   NOR2X0 U366 (.IN1(n205), .IN2(n1193), .QN(n244));
   NOR2X0 U367 (.IN1(n104), .IN2(n95), .QN(n853));
   INVX0 U368 (.INP(n416), .ZN(n1404));
   NOR2X0 U369 (.IN1(n59), .IN2(n48), .QN(n239));
   NOR2X0 U370 (.IN1(n42), .IN2(n62), .QN(n1285));
   NOR2X0 U371 (.IN1(n148), .IN2(n139), .QN(n511));
   NOR2X0 U372 (.IN1(n1285), .IN2(n268), .QN(n1303));
   NOR2X0 U373 (.IN1(n555), .IN2(n500), .QN(n509));
   NOR2X0 U374 (.IN1(n897), .IN2(n842), .QN(n851));
   NOR2X0 U375 (.IN1(n1318), .IN2(n205), .QN(n1345));
   NOR2X0 U376 (.IN1(n1059), .IN2(n868), .QN(n966));
   NOR2X0 U377 (.IN1(n135), .IN2(n150), .QN(n674));
   NOR2X0 U378 (.IN1(n139), .IN2(n147), .QN(n555));
   INVX0 U379 (.INP(n215), .ZN(n49));
   NOR2X0 U380 (.IN1(n159), .IN2(n1406), .QN(n420));
   NOR2X0 U381 (.IN1(n163), .IN2(n1403), .QN(n335));
   NOR2X0 U382 (.IN1(n1405), .IN2(n163), .QN(n480));
   NOR2X0 U383 (.IN1(n842), .IN2(n1069), .QN(n1082));
   INVX0 U384 (.INP(n868), .ZN(n90));
   NOR2X0 U385 (.IN1(n95), .IN2(n103), .QN(n897));
   NOR2X0 U386 (.IN1(n1318), .IN2(n1193), .QN(n1231));
   NOR2X0 U387 (.IN1(n724), .IN2(n526), .QN(n658));
   INVX0 U388 (.INP(n1184), .ZN(n55));
   NOR2X0 U389 (.IN1(n335), .IN2(n280), .QN(n289));
   NOR2X0 U390 (.IN1(n91), .IN2(n108), .QN(n982));
   INVX0 U391 (.INP(n526), .ZN(n134));
   INVX0 U392 (.INP(n306), .ZN(n158));
   NOR2X0 U393 (.IN1(n108), .IN2(n963), .QN(n869));
   NOR2X0 U394 (.IN1(n500), .IN2(n734), .QN(n747));
   NOR2X0 U395 (.IN1(n213), .IN2(n62), .QN(n238));
   NOR2X0 U396 (.IN1(n880), .IN2(n891), .QN(n939));
   NOR2X0 U397 (.IN1(n150), .IN2(n655), .QN(n527));
   NOR2X0 U398 (.IN1(n480), .IN2(n306), .QN(n456));
   NOR2X0 U399 (.IN1(n538), .IN2(n549), .QN(n597));
   NOR2X0 U400 (.IN1(n318), .IN2(n329), .QN(n377));
   INVX0 U401 (.INP(n1280), .ZN(n46));
   NOR2X0 U402 (.IN1(n470), .IN2(n306), .QN(n404));
   INVX0 U403 (.INP(n975), .ZN(n99));
   NOR2X0 U404 (.IN1(n1404), .IN2(n163), .QN(n291));
   INVX0 U405 (.INP(n667), .ZN(n143));
   INVX0 U406 (.INP(n413), .ZN(n167));
   NOR2X0 U407 (.IN1(n280), .IN2(n480), .QN(n493));
   INVX0 U408 (.INP(n1207), .ZN(n56));
   INVX0 U409 (.INP(n1105), .ZN(n84));
   NOR2X0 U410 (.IN1(n1406), .IN2(n401), .QN(n307));
   INVX0 U411 (.INP(n1193), .ZN(n38));
   NOR2X0 U412 (.IN1(n238), .IN2(n1193), .QN(n200));
   INVX0 U413 (.INP(n770), .ZN(n128));
   INVX0 U414 (.INP(n891), .ZN(n98));
   NOR2X0 U415 (.IN1(n238), .IN2(n1262), .QN(n254));
   NOR2X0 U416 (.IN1(n869), .IN2(n1064), .QN(n956));
   INVX0 U417 (.INP(n549), .ZN(n142));
   INVX0 U418 (.INP(n329), .ZN(n166));
   INVX0 U419 (.INP(n273), .ZN(n57));
   NOR2X0 U420 (.IN1(n527), .IN2(n729), .QN(n648));
   INVX0 U421 (.INP(n523), .ZN(n146));
   INVX0 U422 (.INP(n865), .ZN(n102));
   INVX0 U423 (.INP(n1064), .ZN(n83));
   NOR2X0 U424 (.IN1(n869), .IN2(n868), .QN(n959));
   INVX0 U425 (.INP(n1262), .ZN(n34));
   INVX0 U426 (.INP(n729), .ZN(n127));
   INVX0 U427 (.INP(n618), .ZN(n152));
   NOR2X0 U428 (.IN1(n527), .IN2(n526), .QN(n651));
   NOR2X0 U429 (.IN1(n307), .IN2(n306), .QN(n397));
   INVX0 U430 (.INP(n221), .ZN(n33));
   NOR2X0 U431 (.IN1(n880), .IN2(n1065), .QN(n1061));
   NOR2X0 U432 (.IN1(n1202), .IN2(n240), .QN(n195));
   NOR2X0 U433 (.IN1(n538), .IN2(n730), .QN(n726));
   INVX0 U434 (.INP(n550), .ZN(n132));
   INVX0 U435 (.INP(n892), .ZN(n88));
   NOR2X0 U436 (.IN1(n307), .IN2(n475), .QN(n394));
   INVX0 U437 (.INP(n303), .ZN(n1402));
   INVX0 U438 (.INP(n475), .ZN(n151));
   NOR2X0 U439 (.IN1(n95), .IN2(n108), .QN(n1065));
   NOR2X0 U440 (.IN1(n48), .IN2(n62), .QN(n240));
   NOR2X0 U441 (.IN1(n139), .IN2(n150), .QN(n730));
   NOR2X0 U442 (.IN1(n163), .IN2(n1406), .QN(n476));
   INVX0 U443 (.INP(n330), .ZN(n156));
   NOR2X0 U444 (.IN1(n318), .IN2(n476), .QN(n472));
   NOR2X0 U445 (.IN1(n59), .IN2(n62), .QN(n269));
   NOR2X0 U446 (.IN1(n150), .IN2(n147), .QN(n525));
   NOR2X0 U447 (.IN1(n108), .IN2(n103), .QN(n867));
   NOR2X0 U448 (.IN1(n1406), .IN2(n1403), .QN(n305));
   NOR2X0 U449 (.IN1(n65), .IN2(n66), .QN(n172));
   NOR2X0 U450 (.IN1(n110), .IN2(n109), .QN(n1085));
   NOR2X0 U451 (.IN1(n170), .IN2(n169), .QN(n750));
   NOR2X0 U452 (.IN1(n1408), .IN2(n1407), .QN(n598));
   NOR2X0 U453 (.IN1(n15), .IN2(sboxw[22]), .QN(n870));
   NAND2X1 U454 (.IN1(n1127), .IN2(n1128), .QN(n1126));
   INVX0 U455 (.INP(n16), .ZN(n15));
   AO22X1 U456 (.IN1(n15), .IN2(n968), .IN3(n969), .IN4(n16), .Q(n941));
   NAND2X1 U457 (.IN1(sboxw[20]), .IN2(n9), .QN(n954));
   AO22X1 U458 (.IN1(n15), .IN2(n1106), .IN3(n1107), .IN4(n16), .Q(n1088));
   AO22X1 U459 (.IN1(n15), .IN2(n1113), .IN3(n1114), .IN4(n16), .Q(n1086));
   AO22X1 U460 (.IN1(n15), .IN2(n929), .IN3(n930), .IN4(n16), .Q(n901));
   NAND2X1 U461 (.IN1(n15), .IN2(n866), .QN(n855));
   NAND2X1 U462 (.IN1(n918), .IN2(n986), .QN(n980));
   INVX0 U463 (.INP(n934), .ZN(n72));
   INVX0 U464 (.INP(n1061), .ZN(n93));
   AO22X1 U465 (.IN1(n15), .IN2(n911), .IN3(n912), .IN4(n16), .Q(n904));
   NAND2X1 U466 (.IN1(n87), .IN2(n75), .QN(n1154));
   OA222X1 U467 (.IN1(n84), .IN2(n82), .IN3(n15), .IN4(n1162), .IN5(n1163), .IN6(n16), .Q(
          n1161));
   NOR2X0 U468 (.IN1(n106), .IN2(n4), .QN(n302));
   INVX0 U469 (.INP(n5), .ZN(n106));
   NAND2X1 U470 (.IN1(n303), .IN2(n22), .QN(n300));
   NAND2X1 U471 (.IN1(n13), .IN2(n304), .QN(n293));
   NAND2X1 U472 (.IN1(n299), .IN2(n14), .QN(n295));
   NOR2X0 U473 (.IN1(n81), .IN2(n9), .QN(n864));
   INVX0 U474 (.INP(n10), .ZN(n81));
   NAND2X1 U475 (.IN1(n865), .IN2(n71), .QN(n862));
   INVX0 U476 (.INP(n472), .ZN(n161));
   INVX0 U477 (.INP(n882), .ZN(n70));
   OA21X1 U478 (.IN1(n319), .IN2(n158), .IN3(n409), .Q(n450));
   OA21X1 U479 (.IN1(n881), .IN2(n90), .IN3(n971), .Q(n1012));
   INVX0 U480 (.INP(n320), .ZN(n21));
   NAND2X1 U481 (.IN1(n413), .IN2(n319), .QN(n1039));
   NAND2X1 U482 (.IN1(n975), .IN2(n881), .QN(n1136));
   NAND2X1 U483 (.IN1(n155), .IN2(n26), .QN(n1383));
   NAND2X1 U484 (.IN1(n5), .IN2(n622), .QN(n1034));
   NAND2X1 U485 (.IN1(n10), .IN2(n1109), .QN(n1131));
   OA21X1 U486 (.IN1(n896), .IN2(sboxw[18]), .IN3(n78), .Q(n917));
   OA21X1 U487 (.IN1(n334), .IN2(sboxw[2]), .IN3(n29), .Q(n355));
   NAND2X1 U488 (.IN1(n576), .IN2(n678), .QN(n672));
   NAND2X1 U489 (.IN1(n792), .IN2(n793), .QN(n791));
   NAND2X1 U490 (.IN1(sboxw[28]), .IN2(n11), .QN(n646));
   NAND2X1 U491 (.IN1(n667), .IN2(n12), .QN(n742));
   INVX0 U492 (.INP(n726), .ZN(n137));
   OA21X1 U493 (.IN1(n508), .IN2(n509), .IN3(n510), .Q(n507));
   NOR2X0 U494 (.IN1(n13), .IN2(sboxw[6]), .QN(n308));
   NAND2X1 U495 (.IN1(n1030), .IN2(n1031), .QN(n1029));
   NAND2X1 U496 (.IN1(sboxw[4]), .IN2(n4), .QN(n392));
   NAND2X1 U497 (.IN1(n356), .IN2(n424), .QN(n418));
   INVX0 U498 (.INP(n372), .ZN(n23));
   OA21X1 U499 (.IN1(n288), .IN2(n289), .IN3(n290), .Q(n287));
   NOR2X0 U500 (.IN1(n27), .IN2(n5), .QN(n328));
   INVX0 U501 (.INP(n4), .ZN(n27));
   NOR2X0 U502 (.IN1(n76), .IN2(n10), .QN(n890));
   INVX0 U503 (.INP(n9), .ZN(n76));
   NOR2X0 U504 (.IN1(n120), .IN2(n12), .QN(n548));
   INVX0 U505 (.INP(n11), .ZN(n120));
   INVX0 U506 (.INP(n12), .ZN(n125));
   INVX0 U507 (.INP(n6), .ZN(n1412));
   NOR2X0 U508 (.IN1(n1412), .IN2(n7), .QN(n193));
   INVX0 U509 (.INP(n195), .ZN(n36));
   NAND2X1 U510 (.IN1(n8), .IN2(n1359), .QN(n1354));
   NAND2X1 U511 (.IN1(n186), .IN2(n187), .QN(n185));
   OA21X1 U512 (.IN1(n539), .IN2(n134), .IN3(n663), .Q(n704));
   INVX0 U513 (.INP(n7), .ZN(n1415));
   NAND2X1 U514 (.IN1(n667), .IN2(n539), .QN(n801));
   OA21X1 U515 (.IN1(n4), .IN2(n404), .IN3(n405), .Q(n402));
   OA21X1 U516 (.IN1(n9), .IN2(n966), .IN3(n967), .Q(n964));
   NOR2X0 U517 (.IN1(n761), .IN2(n762), .QN(n760));
   OA21X1 U518 (.IN1(n11), .IN2(n658), .IN3(n659), .Q(n656));
   NAND2X1 U519 (.IN1(n519), .IN2(n17), .QN(n515));
   NAND2X1 U520 (.IN1(n523), .IN2(n115), .QN(n520));
   INVX0 U521 (.INP(n540), .ZN(n114));
   NAND2X1 U522 (.IN1(n1262), .IN2(n1409), .QN(n1278));
   OA21X1 U523 (.IN1(n41), .IN2(n1409), .IN3(n1274), .Q(n1310));
   NAND2X1 U524 (.IN1(n194), .IN2(n215), .QN(n211));
   NAND2X1 U525 (.IN1(n443), .IN2(n444), .QN(n429));
   NAND2X1 U526 (.IN1(n1005), .IN2(n1006), .QN(n991));
   NAND2X1 U527 (.IN1(n273), .IN2(n1411), .QN(n1191));
   NOR2X0 U528 (.IN1(n1185), .IN2(n1186), .QN(n1175));
   INVX0 U529 (.INP(n1187), .ZN(n44));
   NAND2X1 U530 (.IN1(n697), .IN2(n698), .QN(n683));
   NOR2X0 U531 (.IN1(n475), .IN2(n476), .QN(n474));
   NOR2X0 U532 (.IN1(n1064), .IN2(n1065), .QN(n1063));
   NAND2X1 U533 (.IN1(n302), .IN2(n163), .QN(n326));
   NAND2X1 U534 (.IN1(n864), .IN2(n95), .QN(n888));
   NOR2X0 U535 (.IN1(n729), .IN2(n730), .QN(n728));
   NAND2X1 U536 (.IN1(n522), .IN2(n139), .QN(n546));
   OA21X1 U537 (.IN1(n554), .IN2(sboxw[26]), .IN3(n2), .Q(n575));
   NOR2X0 U538 (.IN1(n1262), .IN2(n240), .QN(n1330));
   INVX0 U539 (.INP(n262), .ZN(n50));
   NAND2X1 U540 (.IN1(n215), .IN2(n7), .QN(n1341));
   NAND2X1 U541 (.IN1(n1304), .IN2(n1305), .QN(n1290));
   NOR2X0 U542 (.IN1(n5), .IN2(n4), .QN(n319));
   NOR2X0 U543 (.IN1(n10), .IN2(n9), .QN(n881));
   NOR2X0 U544 (.IN1(n12), .IN2(n11), .QN(n539));
   NAND2X1 U545 (.IN1(n6), .IN2(sboxw[12]), .QN(n1259));
   NAND2X1 U546 (.IN1(n12), .IN2(n774), .QN(n796));
   OA21X1 U547 (.IN1(n188), .IN2(sboxw[10]), .IN3(n1), .Q(n1228));
   NOR2X0 U548 (.IN1(n7), .IN2(n6), .QN(n194));
   INVX0 U549 (.INP(n8), .ZN(n64));
   NOR2X0 U550 (.IN1(n64), .IN2(n7), .QN(n206));
   NAND2X1 U551 (.IN1(n7), .IN2(n201), .QN(n198));
   NOR2X0 U552 (.IN1(n64), .IN2(sboxw[14]), .QN(n184));
   NOR2X0 U553 (.IN1(n61), .IN2(sboxw[10]), .QN(n1318));
   NOR2X0 U554 (.IN1(sboxw[11]), .IN2(sboxw[12]), .QN(n250));
   NAND2X1 U555 (.IN1(n868), .IN2(n10), .QN(n914));
   NAND2X1 U556 (.IN1(n306), .IN2(n5), .QN(n352));
   NAND2X1 U557 (.IN1(n842), .IN2(n9), .QN(n924));
   NAND2X1 U558 (.IN1(n280), .IN2(n4), .QN(n362));
   NAND2X1 U559 (.IN1(n500), .IN2(n11), .QN(n582));
   NAND2X1 U560 (.IN1(n335), .IN2(n5), .QN(n322));
   NAND2X1 U561 (.IN1(n897), .IN2(n10), .QN(n884));
   NOR2X0 U562 (.IN1(n60), .IN2(sboxw[10]), .QN(n268));
   NOR2X0 U563 (.IN1(n62), .IN2(sboxw[11]), .QN(n1202));
   NAND2X1 U564 (.IN1(n420), .IN2(n5), .QN(n477));
   NAND2X1 U565 (.IN1(n982), .IN2(n10), .QN(n1066));
   NOR2X0 U566 (.IN1(n105), .IN2(sboxw[18]), .QN(n1059));
   NOR2X0 U567 (.IN1(n108), .IN2(sboxw[19]), .QN(n880));
   NAND2X1 U568 (.IN1(n413), .IN2(n5), .QN(n488));
   NAND2X1 U569 (.IN1(n526), .IN2(n12), .QN(n572));
   NAND2X1 U570 (.IN1(n975), .IN2(n10), .QN(n1077));
   NAND2X1 U571 (.IN1(n555), .IN2(n12), .QN(n542));
   NAND2X1 U572 (.IN1(n674), .IN2(n12), .QN(n731));
   NAND2X1 U573 (.IN1(n470), .IN2(n4), .QN(n457));
   NAND2X1 U574 (.IN1(n1059), .IN2(n9), .QN(n1019));
   NOR2X0 U575 (.IN1(n8), .IN2(sboxw[14]), .QN(n182));
   NOR2X0 U576 (.IN1(n148), .IN2(sboxw[26]), .QN(n500));
   NOR2X0 U577 (.IN1(sboxw[27]), .IN2(sboxw[28]), .QN(n670));
   NOR2X0 U578 (.IN1(n104), .IN2(sboxw[18]), .QN(n842));
   NOR2X0 U579 (.IN1(sboxw[19]), .IN2(sboxw[20]), .QN(n978));
   NOR2X0 U580 (.IN1(n149), .IN2(sboxw[26]), .QN(n724));
   NOR2X0 U581 (.IN1(n150), .IN2(sboxw[27]), .QN(n538));
   NAND2X1 U582 (.IN1(n724), .IN2(n11), .QN(n711));
   NAND2X1 U583 (.IN1(n1105), .IN2(n10), .QN(n1002));
   NAND2X1 U584 (.IN1(n618), .IN2(n5), .QN(n440));
   NOR2X0 U585 (.IN1(n65), .IN2(n8), .QN(n177));
   NAND2X1 U586 (.IN1(n770), .IN2(n12), .QN(n694));
   NAND2X1 U587 (.IN1(n480), .IN2(n4), .QN(n324));
   NAND2X1 U588 (.IN1(n1069), .IN2(n9), .QN(n886));
   NOR2X0 U589 (.IN1(n1404), .IN2(sboxw[2]), .QN(n280));
   NOR2X0 U590 (.IN1(n1405), .IN2(sboxw[2]), .QN(n470));
   NAND2X1 U591 (.IN1(n7), .IN2(n239), .QN(n209));
   OA21X1 U592 (.IN1(n6), .IN2(n34), .IN3(n209), .Q(n1204));
   NAND2X1 U593 (.IN1(n734), .IN2(n11), .QN(n544));
   NAND2X1 U594 (.IN1(n1193), .IN2(n7), .QN(n202));
   NAND2X1 U595 (.IN1(n1285), .IN2(n7), .QN(n1331));
   NOR2X0 U596 (.IN1(n1406), .IN2(sboxw[3]), .QN(n318));
   NOR2X0 U597 (.IN1(sboxw[3]), .IN2(sboxw[4]), .QN(n416));
   INVX0 U598 (.INP(sboxw[10]), .ZN(n48));
   NAND2X1 U599 (.IN1(n6), .IN2(n268), .QN(n1316));
   NAND2X1 U600 (.IN1(n1280), .IN2(n7), .QN(n248));
   NAND2X1 U601 (.IN1(n205), .IN2(n6), .QN(n1205));
   INVX0 U602 (.INP(sboxw[26]), .ZN(n139));
   NOR2X0 U603 (.IN1(sboxw[10]), .IN2(sboxw[12]), .QN(n215));
   INVX0 U604 (.INP(sboxw[2]), .ZN(n163));
   INVX0 U605 (.INP(sboxw[18]), .ZN(n95));
   NOR2X0 U606 (.IN1(n91), .IN2(sboxw[20]), .QN(n868));
   NOR2X0 U607 (.IN1(n62), .IN2(sboxw[10]), .QN(n1184));
   NOR2X0 U608 (.IN1(n135), .IN2(sboxw[28]), .QN(n526));
   NOR2X0 U609 (.IN1(n159), .IN2(sboxw[4]), .QN(n306));
   NAND2X1 U610 (.IN1(sboxw[19]), .IN2(n95), .QN(n963));
   NAND2X1 U611 (.IN1(sboxw[11]), .IN2(n48), .QN(n213));
   NOR2X0 U612 (.IN1(n108), .IN2(sboxw[18]), .QN(n891));
   NAND2X1 U613 (.IN1(sboxw[27]), .IN2(n139), .QN(n655));
   NOR2X0 U614 (.IN1(n150), .IN2(sboxw[26]), .QN(n549));
   NOR2X0 U615 (.IN1(n1406), .IN2(sboxw[2]), .QN(n329));
   NOR2X0 U616 (.IN1(n213), .IN2(sboxw[12]), .QN(n1280));
   NOR2X0 U617 (.IN1(sboxw[18]), .IN2(sboxw[20]), .QN(n975));
   NOR2X0 U618 (.IN1(sboxw[26]), .IN2(sboxw[28]), .QN(n667));
   NOR2X0 U619 (.IN1(sboxw[2]), .IN2(sboxw[4]), .QN(n413));
   INVX0 U620 (.INP(sboxw[12]), .ZN(n62));
   NOR2X0 U621 (.IN1(sboxw[18]), .IN2(sboxw[19]), .QN(n895));
   NOR2X0 U622 (.IN1(sboxw[10]), .IN2(sboxw[11]), .QN(n1207));
   NOR2X0 U623 (.IN1(n42), .IN2(sboxw[12]), .QN(n1193));
   NOR2X0 U624 (.IN1(n963), .IN2(sboxw[20]), .QN(n1105));
   NAND2X1 U625 (.IN1(sboxw[3]), .IN2(n163), .QN(n401));
   NOR2X0 U626 (.IN1(sboxw[26]), .IN2(sboxw[27]), .QN(n553));
   NOR2X0 U627 (.IN1(sboxw[2]), .IN2(sboxw[3]), .QN(n333));
   NOR2X0 U628 (.IN1(n655), .IN2(sboxw[28]), .QN(n770));
   INVX0 U629 (.INP(sboxw[20]), .ZN(n108));
   INVX0 U630 (.INP(sboxw[11]), .ZN(n59));
   INVX0 U631 (.INP(sboxw[28]), .ZN(n150));
   INVX0 U632 (.INP(sboxw[27]), .ZN(n147));
   NOR2X0 U633 (.IN1(n59), .IN2(sboxw[12]), .QN(n273));
   INVX0 U634 (.INP(sboxw[19]), .ZN(n103));
   NOR2X0 U635 (.IN1(n147), .IN2(sboxw[28]), .QN(n523));
   NOR2X0 U636 (.IN1(n103), .IN2(sboxw[20]), .QN(n865));
   NOR2X0 U637 (.IN1(n95), .IN2(sboxw[19]), .QN(n1064));
   NOR2X0 U638 (.IN1(n48), .IN2(sboxw[11]), .QN(n1262));
   NOR2X0 U639 (.IN1(n139), .IN2(sboxw[27]), .QN(n729));
   NOR2X0 U640 (.IN1(n401), .IN2(sboxw[4]), .QN(n618));
   NOR2X0 U641 (.IN1(n48), .IN2(sboxw[12]), .QN(n221));
   NOR2X0 U642 (.IN1(n139), .IN2(sboxw[28]), .QN(n550));
   NOR2X0 U643 (.IN1(n95), .IN2(sboxw[20]), .QN(n892));
   NOR2X0 U644 (.IN1(n66), .IN2(sboxw[14]), .QN(n174));
   INVX0 U645 (.INP(sboxw[4]), .ZN(n1406));
   INVX0 U646 (.INP(sboxw[3]), .ZN(n1403));
   NOR2X0 U647 (.IN1(sboxw[14]), .IN2(sboxw[15]), .QN(n1212));
   NOR2X0 U648 (.IN1(n110), .IN2(sboxw[22]), .QN(n1087));
   NOR2X0 U649 (.IN1(n170), .IN2(sboxw[30]), .QN(n752));
   NOR2X0 U650 (.IN1(n1403), .IN2(sboxw[4]), .QN(n303));
   NOR2X0 U651 (.IN1(sboxw[22]), .IN2(sboxw[23]), .QN(n900));
   NOR2X0 U652 (.IN1(sboxw[30]), .IN2(sboxw[31]), .QN(n558));
   NOR2X0 U653 (.IN1(n163), .IN2(sboxw[3]), .QN(n475));
   NOR2X0 U654 (.IN1(n163), .IN2(sboxw[4]), .QN(n330));
   NOR2X0 U655 (.IN1(n1408), .IN2(sboxw[6]), .QN(n600));
   NOR2X0 U656 (.IN1(sboxw[6]), .IN2(sboxw[7]), .QN(n338));
   NOR2X0 U657 (.IN1(n65), .IN2(sboxw[15]), .QN(n1210));
   NOR2X0 U658 (.IN1(n109), .IN2(sboxw[23]), .QN(n898));
   INVX0 U659 (.INP(sboxw[14]), .ZN(n65));
   INVX0 U660 (.INP(sboxw[22]), .ZN(n109));
   INVX0 U661 (.INP(sboxw[30]), .ZN(n169));
   NOR2X0 U662 (.IN1(n1407), .IN2(sboxw[7]), .QN(n336));
   NOR2X0 U663 (.IN1(n169), .IN2(sboxw[31]), .QN(n556));
   INVX0 U664 (.INP(sboxw[6]), .ZN(n1407));
   INVX0 U665 (.INP(sboxw[15]), .ZN(n66));
   INVX0 U666 (.INP(sboxw[23]), .ZN(n110));
   INVX0 U667 (.INP(sboxw[7]), .ZN(n1408));
   INVX0 U668 (.INP(sboxw[31]), .ZN(n170));
   INVX0 U669 (.INP(sboxw[21]), .ZN(n16));
   NBUFFX4 U670 (.INP(sboxw[1]), .Z(n5));
   NBUFFX4 U671 (.INP(sboxw[17]), .Z(n10));
   NBUFFX4 U672 (.INP(sboxw[25]), .Z(n12));
   INVX0 U673 (.INP(n219), .ZN(n1));
   INVX0 U674 (.INP(n219), .ZN(n1414));
   NOR2X0 U675 (.IN1(n1415), .IN2(n6), .QN(n219));
   INVX0 U676 (.INP(n522), .ZN(n2));
   INVX0 U677 (.INP(n522), .ZN(n122));
   NOR2X0 U930 (.IN1(n125), .IN2(n11), .QN(n522));
   NOR2X0 U931 (.IN1(n17), .IN2(n12), .QN(n501));
   NOR2X0 U1077 (.IN1(n169), .IN2(n17), .QN(n638));
   NOR2X0 U1086 (.IN1(n17), .IN2(sboxw[30]), .QN(n530));
   AO221X1 U1110 (.IN1(n3), .IN2(n672), .IN3(n673), .IN4(n17), .IN5(n116), .Q(n671));
   INVX0 U1203 (.INP(n864), .ZN(n78));
   INVX0 U1209 (.INP(n302), .ZN(n29));
   INVX0 U1251 (.INP(n592), .ZN(n116));
   INVX0 U1434 (.INP(n14), .ZN(n13));
   NOR2X0 U1435 (.IN1(n14), .IN2(n5), .QN(n281));
   NOR2X0 U1436 (.IN1(n1407), .IN2(n14), .QN(n384));
   NOR2X0 U1437 (.IN1(n14), .IN2(sboxw[6]), .QN(n310));
   NAND2X0 U1438 (.IN1(n3), .IN2(n524), .QN(n513));
   NAND2X0 U1439 (.IN1(n3), .IN2(n763), .QN(n758));
   NOR2X0 U1440 (.IN1(n3), .IN2(sboxw[30]), .QN(n528));
   NOR2X0 U1441 (.IN1(n169), .IN2(n3), .QN(n640));
   INVX0 U1442 (.INP(sboxw[5]), .ZN(n14));
   NAND2X0 U1443 (.IN1(n861), .IN2(n16), .QN(n857));
   NOR2X0 U1444 (.IN1(n109), .IN2(n16), .QN(n946));
   NOR2X0 U1445 (.IN1(n16), .IN2(sboxw[22]), .QN(n872));
   NOR2X0 U1446 (.IN1(n16), .IN2(n10), .QN(n843));
   INVX0 U1447 (.INP(sboxw[29]), .ZN(n17));
endmodule

module aes_decipher_block_test_1 (clk, reset_n, next, keylen, round, round_key, block, 
       new_block, ready, test_si, test_so, test_se);
input clk, reset_n, next, keylen, test_si, test_se;
input [127:0] round_key;
input [127:0] block;
output ready, test_so;
output [3:0] round;
output [127:0] new_block;
wire n158, n159, n164, n166, n167, n169, n170, n171, n172, n173, n177, n180, n182, n184, 
       n185, n186, n187, n188, n190, n193, n195, n197, n199, n200, n201, n202, n203, n204
       , n205, n209, n211, n213, n215, n216, n217, n218, n219, n222, n225, n227, n229, 
       n230, n231, n232, n233, n234, n237, n239, n241, n243, n244, n245, n246, n253, n256
       , n258, n260, n261, n262, n263, n264, n265, n270, n272, n274, n275, n276, n277, 
       n278, n280, n284, n286, n288, n289, n290, n291, n292, n296, n298, n300, n302, n303
       , n304, n305, n306, n307, n313, n315, n317, n318, n319, n321, n322, n323, n326, 
       n328, n330, n332, n333, n334, n335, n464, n465, n466, n467, n468, n469, n470, n471
       , n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
       n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498
       , n499, n501, n502, n503, n504, n505, n507, n508, n509, n510, n511, n512, n513, 
       n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n526, n527, n528
       , n529, n530, n531, n532, n533, n534, n535, n536, n537, n539, n540, n541, n542, 
       n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557
       , n558, n559, n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571, 
       n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n585, n586
       , n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n600, 
       n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614
       , n615, n616, n617, n618, n620, n621, n622, n623, n624, n626, n627, n628, n629, 
       n630, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644
       , n645, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
       n659, n660, n661, n662, n663, n665, n666, n667, n668, n669, n670, n671, n672, n673
       , n674, n675, n676, n677, n678, n680, n681, n682, n683, n684, n685, n686, n687, 
       n688, n689, n690, n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702
       , n703, n704, n705, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, 
       n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n728, n729, n730, n731
       , n732, n733, n734, n735, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
       n746, n747, n748, n749, n750, n751, n752, n754, n755, n756, n757, n758, n759, n760
       , n761, n762, n763, n764, n765, n766, n767, n769, n770, n771, n772, n773, n774, 
       n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n787, n788, n789, n790
       , n791, n792, n793, n794, n795, n796, n797, n798, n799, n801, n802, n803, n804, 
       n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n817, n818, n819
       , n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n835, 
       n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849
       , n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, 
       n864, n865, n866, n867, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878
       , n879, n880, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, 
       n893, n894, n895, n896, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907
       , n908, n909, n910, n911, n912, n913, n915, n916, n917, n918, n919, n920, n921, 
       n922, n923, n924, n925, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936
       , n937, n938, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
       n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964
       , n965, n966, n967, n968, n969, n970, n972, n973, n974, n975, n976, n977, n978, 
       n980, n981, n982, n983, n984, n986, n987, n988, n989, n990, n991, n992, n993, n994
       , n995, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, 
       n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020
       , n1021, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
       n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045
       , n1046, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, 
       n1058, n1059, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070
       , n1071, n1072, n1073, n1074, n1075, n1077, n1078, n1079, n1080, n1082, n1083, 
       n1084, n1085, n1086, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098
       , n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, 
       n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124
       , n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1134, n1135, n1136, n1137, 
       n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1147, n1148, n1149, n1150
       , n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
       n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1170, n1171, n1172, n1173, n1174
       , n1175, n1176, n1177, n1178, n1179, n1181, n1182, n1183, n1184, n1185, n1186, 
       n1187, n1188, n1189, n1190, n1191, n1194, n1195, n1196, n1197, n1198, n1199, n1200
       , n1201, n1202, n1204, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
       n1214, n1215, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228
       , n1229, n1230, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
       n1241, n1242, n1243, n1244, n1245, n1246, n1249, n1250, n1251, n1252, n1253, n1254
       , n1255, n1256, n1257, n1258, n1259, n1260, n1264, n1265, n1266, n1267, n1268, 
       n1269, n1270, n1271, n1272, n1273, n1277, n1278, n1279, n1280, n1281, n1282, n1283
       , n1284, n1285, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1298, 
       n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1311
       , n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
       n1323, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335
       , n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
       n1347, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359
       , n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1373, n1374, 
       n1375, n1376, n1378, n1379, n1380, n1381, n1383, n1384, n1385, n1386, n1387, n1388
       , n1389, n1393, n1394, n1395, n1396, n1397, n1398, n1400, n1401, n1402, n1403, 
       n1404, n1405, n1406, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1417
       , n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
       n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1441
       , n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1451, n1452, n1453, 
       n1454, n1455, n1456, n1457, n1458, n1459, n1461, n1462, n1463, n1464, n1465, n1466
       , n1467, n1468, n1469, n1471, n1472, n1473, n1474, n1475, n1476, n1478, n1479, 
       n1480, n1481, n1482, n1483, n1484, n1485, n1487, n1488, n1489, n1490, n1491, n1492
       , n1493, n1494, n1495, n1496, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
       n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516
       , n1517, n1518, n1519, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1529, 
       n1531, n1532, n1533, n1534, n1535, n1536, n1540, n1541, n1542, n1543, n1544, n1545
       , n1546, n1547, n1550, n1551, n1552, n1553, n1554, n1555, n1557, n1558, n1559, 
       n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572
       , n1573, n1574, n1575, n1576, n1577, n1578, n1580, n1581, n1582, n1583, n1584, 
       n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1596, n1597, n1598
       , n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1607, n1608, n1609, n1610, 
       n1611, n1612, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1624, n1625, n1626
       , n1627, n1628, n1629, n1630, n1631, n1633, n1635, n1636, n1637, n1638, n1639, 
       n1640, n1641, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1652, n1653
       , n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1662, n1663, n1664, n1665, 
       n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1675, n1676, n1677, n1678
       , n1679, n1680, n1681, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, 
       n1694, n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1704, n1705, n1706, n1707
       , n1708, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1720, 
       n1721, n1722, n1723, n1724, n1725, n1727, n1728, n1729, n1730, n1731, n1732, n1733
       , n1734, n1735, n1736, n1737, n1739, n1740, n1741, n1742, n1743, n1745, n1746, 
       n1747, n1748, n1749, n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1758, n1759
       , n1761, n1762, n1763, n1765, n1766, n1767, n1768, n1769, n1773, n1774, n1775, 
       n1776, n1777, n1778, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1789
       , n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, 
       n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1810, n1811, n1812, n1813, n1814
       , n1815, n1816, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1827, 
       n1828, n1829, n1830, n1831, n1832, n1833, n1835, n1836, n1837, n1838, n1839, n1840
       , n1841, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1853, 
       n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1864, n1865, n1866, n1867, n1868
       , n1869, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
       n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1893, n1894, n1895, n1896
       , n1897, n1898, n1899, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1913, 
       n1914, n1915, n1916, n1917, n1918, n1920, n1921, n1922, n1923, n1924, n1925, n1927
       , n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1936, n1937, n1938, n1939, 
       n1940, n1941, n1942, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952
       , n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1963, n1964, n1965, 
       n1966, n1967, n1968, n1969, n1971, n1972, n1973, n1974, n1975, n1976, n1978, n1979
       , n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1989, n1990, n1991, 
       n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003
       , n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, 
       n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026
       , n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
       n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049
       , n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
       n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072
       , n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
       n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095
       , n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, 
       n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118
       , n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
       n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141
       , n2142, n1, n2, n3, n4, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151
       , n152, n153, n154, n155, n156, n157, n160, n161, n162, n163, n165, n168, n174, 
       n175, n176, n178, n179, n181, n183, n189, n191, n192, n194, n196, n198, n206, n207
       , n208, n210, n212, n214, n220, n221, n223, n224, n226, n228, n235, n236, n238, 
       n240, n242, n247, n248, n249, n250, n251, n252, n254, n255, n257, n259, n266, n267
       , n268, n269, n271, n273, n279, n281, n282, n283, n285, n287, n293, n294, n295, 
       n297, n299, n301, n308, n309, n310, n311, n312, n314, n316, n320, n324, n325, n327
       , n329, n331, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
       n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360
       , n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
       n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387
       , n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
       n401, n402, n403, n404, n405, n406, n407, n408, n409, n434, n435, n436, n437, n438
       , n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
       n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n500, n506
       , n525, n538, n553, n567, n584, n599, n619, n625, n631, n646, n664, n679, n697, 
       n706, n727, n736, n753, n768, n785, n786, n800, n816, n832, n833, n834, n850, n868
       , n881, n897, n914, n926, n939, n971, n979, n985, n996, n1008, n1022, n1033, n1047
       , n1060, n1076, n1081, n1087, n1088, n1089, n1099, n1100, n1112, n1125, n1133, 
       n1146, n1169, n1180, n1192, n1193, n1203, n1205, n1216, n1217, n1218, n1231, n1247
       , n1248, n1261, n1262, n1263, n1274, n1275, n1276, n1286, n1287, n1288, n1297, 
       n1310, n1324, n1348, n1360, n1370, n1371, n1372, n1377, n1382, n1390, n1391, n1392
       , n1399, n1407, n1416, n1440, n1450, n1460, n1470, n1477, n1486, n1497, n1520, 
       n1528, n1530, n1537, n1538, n1539, n1548, n1549, n1556, n1568, n1579, n1594, n1595
       , n1606, n1613, n1614, n1615, n1623, n1632, n1634, n1642, n1651, n1661, n1674, 
       n1682, n1691, n1692, n1693, n1696, n1703, n1709, n1719, n1726, n1738, n1744, n1752
       , n1760, n1764, n1770, n1771, n1772, n1779, n1788, n1801, n1809, n1817, n1826, 
       n1834, n1842, n1852, n1861, n1862, n1863, n1870, n1871, n1872, n1883, n1892, n1900
       , n1901, n1902, n1910, n1911, n1912, n1919, n1926, n1935, n1943, n1953, n1962, 
       n1970, n1977, n1988, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151
       , n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
       n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174
       , n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, 
       n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197
       , n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, 
       n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220
       , n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2232, 
       n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244
       , n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, 
       n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267
       ;
wire [31:0] tmp_sboxw;
wire [31:0] new_sboxw;
wire [1:0] sword_ctr_reg;
wire [1:0] dec_ctrl_reg;
   assign test_so = n204;
   SDFFARX1 \sword_ctr_reg_reg[0]  (.D(n2142), .SI(n2232), .SE(test_se), .CLK(clk), .RSTB(
          n1133), .Q(sword_ctr_reg[0]), .QN(n205));
   SDFFARX1 \sword_ctr_reg_reg[1]  (.D(n2141), .SI(sword_ctr_reg[0]), .SE(test_se), .CLK(
          clk), .RSTB(n1089), .Q(sword_ctr_reg[1]), .QN(n204));
   SDFFARX1 \round_ctr_reg_reg[1]  (.D(n2137), .SI(n2234), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(round[1]), .QN(n203));
   SDFFARX1 \round_ctr_reg_reg[2]  (.D(n2136), .SI(n203), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(round[2]), .QN(n2233));
   SDFFARX1 \round_ctr_reg_reg[3]  (.D(n2135), .SI(n2233), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(round[3]), .QN(n2232));
   SDFFASX1 ready_reg_reg (.D(n2134), .SI(dec_ctrl_reg[1]), .SE(test_se), .CLK(clk), .SETB(
          n1203), .Q(ready), .QN(n2235));
   SDFFARX1 \block_w0_reg_reg[0]  (.D(n2133), .SI(test_si), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(new_block[96]), .QN(n335));
   SDFFARX1 \block_w3_reg_reg[1]  (.D(n2131), .SI(new_block[0]), .SE(test_se), .CLK(clk), .
          RSTB(n1089), .Q(new_block[1]), .QN(n201));
   SDFFARX1 \block_w0_reg_reg[31]  (.D(n2006), .SI(n2261), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(new_block[127]), .QN(n2260));
   SDFFARX1 \block_w3_reg_reg[0]  (.D(n2132), .SI(n2244), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[0]), .QN(n202));
   SDFFARX1 \block_w3_reg_reg[24]  (.D(n2108), .SI(new_block[23]), .SE(test_se), .CLK(clk)
          , .RSTB(n1099), .Q(new_block[24]), .QN(n2243));
   SDFFARX1 \block_w3_reg_reg[26]  (.D(n2106), .SI(n2242), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[26]), .QN(n2241));
   SDFFARX1 \block_w3_reg_reg[27]  (.D(n2105), .SI(n2241), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[27]), .QN(n2240));
   SDFFARX1 \block_w0_reg_reg[23]  (.D(n2014), .SI(new_block[118]), .SE(test_se), .CLK(clk)
          , .RSTB(n1099), .Q(new_block[119]), .QN(n296));
   SDFFARX1 \block_w2_reg_reg[15]  (.D(n2085), .SI(new_block[46]), .SE(test_se), .CLK(clk)
          , .RSTB(n1099), .Q(new_block[47]), .QN(n222));
   SDFFARX1 \block_w3_reg_reg[16]  (.D(n2116), .SI(n177), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[16]), .QN(n173));
   SDFFARX1 \block_w2_reg_reg[3]  (.D(n2097), .SI(new_block[34]), .SE(test_se), .CLK(clk)
          , .RSTB(n1099), .Q(new_block[35]), .QN(n243));
   SDFFARX1 \block_w3_reg_reg[19]  (.D(n2113), .SI(new_block[18]), .SE(test_se), .CLK(clk)
          , .RSTB(n1099), .Q(new_block[19]), .QN(n170));
   SDFFARX1 \block_w1_reg_reg[9]  (.D(n2059), .SI(new_block[72]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[73]), .QN(n277));
   SDFFARX1 \block_w3_reg_reg[10]  (.D(n2122), .SI(new_block[9]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[10]), .QN(n186));
   SDFFARX1 \block_w3_reg_reg[3]  (.D(n2129), .SI(new_block[2]), .SE(test_se), .CLK(clk), .
          RSTB(n1100), .Q(new_block[3]), .QN(n199));
   SDFFARX1 \block_w3_reg_reg[15]  (.D(n2117), .SI(new_block[14]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[15]), .QN(n177));
   SDFFARX1 \block_w1_reg_reg[10]  (.D(n2058), .SI(new_block[73]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[74]), .QN(n276));
   SDFFARX1 \block_w2_reg_reg[19]  (.D(n2081), .SI(new_block[50]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[51]), .QN(n216));
   SDFFARX1 \block_w3_reg_reg[20]  (.D(n2112), .SI(new_block[19]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[20]), .QN(n169));
   SDFFARX1 \block_w2_reg_reg[6]  (.D(n2094), .SI(new_block[37]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[38]), .QN(n237));
   SDFFARX1 \block_w2_reg_reg[30]  (.D(n2070), .SI(n2246), .SE(test_se), .CLK(clk), .RSTB(
          n1100), .Q(new_block[62]), .QN(n2245));
   SDFFARX1 \block_w1_reg_reg[7]  (.D(n2061), .SI(new_block[70]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[71]), .QN(n280));
   SDFFARX1 \block_w3_reg_reg[8]  (.D(n2124), .SI(n190), .SE(test_se), .CLK(clk), .RSTB(
          n1112), .Q(new_block[8]), .QN(n188));
   SDFFARX1 \block_w0_reg_reg[17]  (.D(n2020), .SI(new_block[112]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[113]), .QN(n305));
   SDFFARX1 \block_w1_reg_reg[19]  (.D(n2049), .SI(new_block[82]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[83]), .QN(n261));
   SDFFARX1 \block_w3_reg_reg[11]  (.D(n2121), .SI(new_block[10]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[11]), .QN(n185));
   SDFFARX1 \block_w3_reg_reg[4]  (.D(n2128), .SI(new_block[3]), .SE(test_se), .CLK(clk), .
          RSTB(n1112), .Q(new_block[4]), .QN(n197));
   SDFFARX1 \block_w3_reg_reg[7]  (.D(n2125), .SI(new_block[6]), .SE(test_se), .CLK(clk), .
          RSTB(n1112), .Q(new_block[7]), .QN(n190));
   SDFFARX1 \block_w2_reg_reg[1]  (.D(n2099), .SI(new_block[32]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[33]), .QN(n245));
   SDFFARX1 \block_w3_reg_reg[17]  (.D(n2115), .SI(new_block[16]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[17]), .QN(n172));
   SDFFARX1 \block_w1_reg_reg[5]  (.D(n2063), .SI(new_block[68]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[69]), .QN(n286));
   SDFFARX1 \block_w0_reg_reg[6]  (.D(n2031), .SI(new_block[101]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[102]), .QN(n326));
   SDFFARX1 \block_w0_reg_reg[30]  (.D(n2007), .SI(n2262), .SE(test_se), .CLK(clk), .RSTB(
          n1125), .Q(new_block[126]), .QN(n2261));
   SDFFARX1 \block_w1_reg_reg[22]  (.D(n2046), .SI(new_block[85]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[86]), .QN(n256));
   SDFFARX1 \block_w3_reg_reg[13]  (.D(n2119), .SI(new_block[12]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[13]), .QN(n182));
   SDFFARX1 \block_w1_reg_reg[3]  (.D(n2065), .SI(new_block[66]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[67]), .QN(n289));
   SDFFARX1 \block_w1_reg_reg[20]  (.D(n2048), .SI(new_block[83]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[84]), .QN(n260));
   SDFFARX1 \block_w2_reg_reg[22]  (.D(n2078), .SI(new_block[53]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[54]), .QN(n211));
   SDFFARX1 \block_w1_reg_reg[4]  (.D(n2064), .SI(new_block[67]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[68]), .QN(n288));
   SDFFARX1 \block_w0_reg_reg[5]  (.D(n2032), .SI(new_block[100]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[101]), .QN(n328));
   SDFFARX1 \block_w1_reg_reg[21]  (.D(n2047), .SI(new_block[84]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[85]), .QN(n258));
   SDFFARX1 \block_w0_reg_reg[15]  (.D(n2022), .SI(new_block[110]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[111]), .QN(n307));
   SDFFARX1 \block_w3_reg_reg[2]  (.D(n2130), .SI(new_block[1]), .SE(test_se), .CLK(clk), .
          RSTB(n1133), .Q(new_block[2]), .QN(n200));
   SDFFARX1 \block_w0_reg_reg[16]  (.D(n2021), .SI(n307), .SE(test_se), .CLK(clk), .RSTB(
          n1133), .Q(new_block[112]), .QN(n306));
   SDFFARX1 \block_w1_reg_reg[18]  (.D(n2050), .SI(new_block[81]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[82]), .QN(n262));
   SDFFARX1 \block_w1_reg_reg[27]  (.D(n2041), .SI(n2257), .SE(test_se), .CLK(clk), .RSTB(
          n1133), .Q(new_block[91]), .QN(n2256));
   SDFFARX1 \block_w0_reg_reg[7]  (.D(n2030), .SI(new_block[102]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[103]), .QN(n323));
   SDFFARX1 \block_w1_reg_reg[17]  (.D(n2051), .SI(new_block[80]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[81]), .QN(n263));
   SDFFARX1 \block_w3_reg_reg[9]  (.D(n2123), .SI(new_block[8]), .SE(test_se), .CLK(clk), .
          RSTB(n1146), .Q(new_block[9]), .QN(n187));
   SDFFARX1 \block_w1_reg_reg[11]  (.D(n2057), .SI(new_block[74]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[75]), .QN(n275));
   SDFFARX1 \block_w3_reg_reg[14]  (.D(n2118), .SI(new_block[13]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[14]), .QN(n180));
   SDFFARX1 \block_w0_reg_reg[3]  (.D(n2034), .SI(new_block[98]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[99]), .QN(n332));
   SDFFARX1 \block_w3_reg_reg[5]  (.D(n2127), .SI(new_block[4]), .SE(test_se), .CLK(clk), .
          RSTB(n1146), .Q(new_block[5]), .QN(n195));
   SDFFARX1 \block_w2_reg_reg[0]  (.D(n2100), .SI(n2252), .SE(test_se), .CLK(clk), .RSTB(
          n1146), .Q(new_block[32]), .QN(n246));
   SDFFARX1 \block_w3_reg_reg[18]  (.D(n2114), .SI(new_block[17]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[18]), .QN(n171));
   SDFFARX1 \block_w1_reg_reg[6]  (.D(n2062), .SI(new_block[69]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[70]), .QN(n284));
   SDFFARX1 \block_w2_reg_reg[21]  (.D(n2079), .SI(new_block[52]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[53]), .QN(n213));
   SDFFARX1 \block_w2_reg_reg[11]  (.D(n2089), .SI(new_block[42]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[43]), .QN(n230));
   SDFFARX1 \block_w3_reg_reg[22]  (.D(n2110), .SI(new_block[21]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[22]), .QN(n166));
   SDFFARX1 \block_w2_reg_reg[2]  (.D(n2098), .SI(new_block[33]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[34]), .QN(n244));
   SDFFARX1 \block_w3_reg_reg[21]  (.D(n2111), .SI(new_block[20]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[21]), .QN(n167));
   SDFFARX1 \block_w1_reg_reg[8]  (.D(n2060), .SI(new_block[71]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[72]), .QN(n278));
   SDFFARX1 \block_w2_reg_reg[7]  (.D(n2093), .SI(new_block[38]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[39]), .QN(n234));
   SDFFARX1 \block_w1_reg_reg[1]  (.D(n2067), .SI(new_block[64]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[65]), .QN(n291));
   SDFFARX1 \block_w3_reg_reg[12]  (.D(n2120), .SI(new_block[11]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[12]), .QN(n184));
   SDFFARX1 \block_w3_reg_reg[31]  (.D(n2101), .SI(n2237), .SE(test_se), .CLK(clk), .RSTB(
          n1169), .Q(new_block[31]), .QN(n2236));
   SDFFARX1 \block_w0_reg_reg[18]  (.D(n2019), .SI(new_block[113]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[114]), .QN(n304));
   SDFFARX1 \block_w0_reg_reg[27]  (.D(n2010), .SI(n2265), .SE(test_se), .CLK(clk), .RSTB(
          n1180), .Q(new_block[123]), .QN(n2264));
   SDFFARX1 \block_w3_reg_reg[6]  (.D(n2126), .SI(new_block[5]), .SE(test_se), .CLK(clk), .
          RSTB(n1180), .Q(new_block[6]), .QN(n193));
   SDFFARX1 \block_w1_reg_reg[14]  (.D(n2054), .SI(new_block[77]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[78]), .QN(n270));
   SDFFARX1 \block_w1_reg_reg[24]  (.D(n2044), .SI(n253), .SE(test_se), .CLK(clk), .RSTB(
          n1180), .Q(new_block[88]), .QN(n2259));
   SDFFARX1 \block_w1_reg_reg[26]  (.D(n2042), .SI(n2258), .SE(test_se), .CLK(clk), .RSTB(
          n1180), .Q(new_block[90]), .QN(n2257));
   SDFFARX1 \block_w2_reg_reg[18]  (.D(n2082), .SI(new_block[49]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[50]), .QN(n217));
   SDFFARX1 \block_w2_reg_reg[26]  (.D(n2074), .SI(n2250), .SE(test_se), .CLK(clk), .RSTB(
          n1180), .Q(new_block[58]), .QN(n2249));
   SDFFARX1 \block_w3_reg_reg[23]  (.D(n2109), .SI(new_block[22]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[23]), .QN(n164));
   SDFFARX1 \block_w1_reg_reg[15]  (.D(n2053), .SI(new_block[78]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[79]), .QN(n265));
   SDFFARX1 \block_w2_reg_reg[17]  (.D(n2083), .SI(new_block[48]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[49]), .QN(n218));
   SDFFARX1 \block_w0_reg_reg[28]  (.D(n2009), .SI(n2264), .SE(test_se), .CLK(clk), .RSTB(
          n1192), .Q(new_block[124]), .QN(n2263));
   SDFFARX1 \block_w1_reg_reg[23]  (.D(n2045), .SI(new_block[86]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[87]), .QN(n253));
   SDFFARX1 \block_w1_reg_reg[31]  (.D(n2037), .SI(n2253), .SE(test_se), .CLK(clk), .RSTB(
          n1192), .Q(new_block[95]), .QN(n2252));
   SDFFARX1 \block_w2_reg_reg[23]  (.D(n2077), .SI(new_block[54]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[55]), .QN(n209));
   SDFFARX1 \block_w2_reg_reg[31]  (.D(n2069), .SI(n2245), .SE(test_se), .CLK(clk), .RSTB(
          n1192), .Q(new_block[63]), .QN(n2244));
   SDFFARX1 \block_w0_reg_reg[1]  (.D(n2036), .SI(new_block[96]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[97]), .QN(n334));
   SDFFARX1 \block_w2_reg_reg[9]  (.D(n2091), .SI(new_block[40]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[41]), .QN(n232));
   SDFFARX1 \block_w2_reg_reg[25]  (.D(n2075), .SI(n2251), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[57]), .QN(n2250));
   SDFFARX1 \block_w0_reg_reg[9]  (.D(n2028), .SI(new_block[104]), .SE(test_se), .CLK(clk)
          , .RSTB(n1193), .Q(new_block[105]), .QN(n321));
   SDFFARX1 \block_w0_reg_reg[25]  (.D(n2012), .SI(n2267), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[121]), .QN(n2266));
   SDFFARX1 \block_w0_reg_reg[26]  (.D(n2011), .SI(n2266), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[122]), .QN(n2265));
   SDFFARX1 \block_w0_reg_reg[29]  (.D(n2008), .SI(n2263), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[125]), .QN(n2262));
   SDFFARX1 \block_w2_reg_reg[8]  (.D(n2092), .SI(n234), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[40]), .QN(n233));
   SDFFARX1 \block_w2_reg_reg[24]  (.D(n2076), .SI(new_block[55]), .SE(test_se), .CLK(clk)
          , .RSTB(n1193), .Q(new_block[56]), .QN(n2251));
   SDFFARX1 \block_w1_reg_reg[0]  (.D(n2068), .SI(n2260), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[64]), .QN(n292));
   SDFFARX1 \block_w2_reg_reg[16]  (.D(n2084), .SI(new_block[47]), .SE(test_se), .CLK(clk)
          , .RSTB(n1193), .Q(new_block[48]), .QN(n219));
   SDFFARX1 \block_w0_reg_reg[8]  (.D(n2029), .SI(n323), .SE(test_se), .CLK(clk), .RSTB(
          n1193), .Q(new_block[104]), .QN(n322));
   SDFFARX1 \block_w0_reg_reg[24]  (.D(n2013), .SI(new_block[119]), .SE(test_se), .CLK(clk)
          , .RSTB(n1193), .Q(new_block[120]), .QN(n2267));
   SDFFARX1 \block_w0_reg_reg[10]  (.D(n2027), .SI(new_block[105]), .SE(test_se), .CLK(clk)
          , .RSTB(n1193), .Q(new_block[106]), .QN(n319));
   SDFFARX1 \block_w1_reg_reg[16]  (.D(n2052), .SI(n265), .SE(test_se), .CLK(clk), .RSTB(
          n1203), .Q(new_block[80]), .QN(n264));
   SDFFARX1 \block_w0_reg_reg[2]  (.D(n2035), .SI(new_block[97]), .SE(test_se), .CLK(clk)
          , .RSTB(n1203), .Q(new_block[98]), .QN(n333));
   SDFFARX1 \block_w2_reg_reg[10]  (.D(n2090), .SI(new_block[41]), .SE(test_se), .CLK(clk)
          , .RSTB(n1203), .Q(new_block[42]), .QN(n231));
   SDFFARX1 \block_w1_reg_reg[2]  (.D(n2066), .SI(new_block[65]), .SE(test_se), .CLK(clk)
          , .RSTB(n1089), .Q(new_block[66]), .QN(n290));
   AO221X1 U575 (.IN1(new_block[9]), .IN2(n452), .IN3(new_block[41]), .IN4(n456), .IN5(
          n464), .Q(tmp_sboxw[9]));
   AO22X1 U576 (.IN1(new_block[105]), .IN2(n454), .IN3(new_block[73]), .IN4(n450), .Q(n464)
          );
   AO221X1 U577 (.IN1(new_block[8]), .IN2(n451), .IN3(new_block[40]), .IN4(n456), .IN5(
          n465), .Q(tmp_sboxw[8]));
   AO22X1 U578 (.IN1(new_block[104]), .IN2(n453), .IN3(new_block[72]), .IN4(n450), .Q(n465)
          );
   AO221X1 U579 (.IN1(new_block[7]), .IN2(n452), .IN3(new_block[39]), .IN4(n456), .IN5(
          n466), .Q(tmp_sboxw[7]));
   AO22X1 U580 (.IN1(new_block[103]), .IN2(n453), .IN3(new_block[71]), .IN4(n450), .Q(n466)
          );
   AO221X1 U581 (.IN1(new_block[6]), .IN2(n451), .IN3(new_block[38]), .IN4(n456), .IN5(
          n467), .Q(tmp_sboxw[6]));
   AO22X1 U582 (.IN1(new_block[102]), .IN2(n454), .IN3(new_block[70]), .IN4(n450), .Q(n467)
          );
   AO221X1 U583 (.IN1(new_block[5]), .IN2(n452), .IN3(new_block[37]), .IN4(n456), .IN5(
          n468), .Q(tmp_sboxw[5]));
   AO22X1 U584 (.IN1(new_block[101]), .IN2(n453), .IN3(new_block[69]), .IN4(n450), .Q(n468)
          );
   AO221X1 U585 (.IN1(new_block[4]), .IN2(n451), .IN3(new_block[36]), .IN4(n456), .IN5(
          n469), .Q(tmp_sboxw[4]));
   AO22X1 U586 (.IN1(new_block[100]), .IN2(n454), .IN3(new_block[68]), .IN4(n450), .Q(n469)
          );
   AO221X1 U587 (.IN1(new_block[3]), .IN2(n452), .IN3(new_block[35]), .IN4(n456), .IN5(
          n470), .Q(tmp_sboxw[3]));
   AO22X1 U588 (.IN1(new_block[99]), .IN2(n454), .IN3(new_block[67]), .IN4(n450), .Q(n470)
          );
   AO221X1 U589 (.IN1(new_block[31]), .IN2(n451), .IN3(new_block[63]), .IN4(n456), .IN5(
          n471), .Q(tmp_sboxw[31]));
   AO22X1 U590 (.IN1(new_block[127]), .IN2(n454), .IN3(new_block[95]), .IN4(n450), .Q(n471)
          );
   AO221X1 U591 (.IN1(new_block[30]), .IN2(n452), .IN3(new_block[62]), .IN4(n455), .IN5(
          n472), .Q(tmp_sboxw[30]));
   AO221X1 U593 (.IN1(new_block[2]), .IN2(n452), .IN3(new_block[34]), .IN4(n456), .IN5(
          n473), .Q(tmp_sboxw[2]));
   AO221X1 U595 (.IN1(new_block[29]), .IN2(n452), .IN3(new_block[61]), .IN4(n456), .IN5(
          n474), .Q(tmp_sboxw[29]));
   AO221X1 U597 (.IN1(new_block[28]), .IN2(n452), .IN3(new_block[60]), .IN4(n455), .IN5(
          n475), .Q(tmp_sboxw[28]));
   AO221X1 U599 (.IN1(new_block[27]), .IN2(n452), .IN3(new_block[59]), .IN4(n455), .IN5(
          n476), .Q(tmp_sboxw[27]));
   AO221X1 U601 (.IN1(new_block[26]), .IN2(n452), .IN3(new_block[58]), .IN4(n456), .IN5(
          n477), .Q(tmp_sboxw[26]));
   AO221X1 U603 (.IN1(new_block[25]), .IN2(n452), .IN3(new_block[57]), .IN4(n456), .IN5(
          n478), .Q(tmp_sboxw[25]));
   AO221X1 U605 (.IN1(new_block[24]), .IN2(n452), .IN3(new_block[56]), .IN4(n456), .IN5(
          n479), .Q(tmp_sboxw[24]));
   AO221X1 U607 (.IN1(new_block[23]), .IN2(n452), .IN3(new_block[55]), .IN4(n456), .IN5(
          n480), .Q(tmp_sboxw[23]));
   AO221X1 U609 (.IN1(new_block[22]), .IN2(n452), .IN3(new_block[54]), .IN4(n456), .IN5(
          n481), .Q(tmp_sboxw[22]));
   AO221X1 U611 (.IN1(new_block[21]), .IN2(n452), .IN3(new_block[53]), .IN4(n455), .IN5(
          n482), .Q(tmp_sboxw[21]));
   AO221X1 U613 (.IN1(new_block[20]), .IN2(n452), .IN3(new_block[52]), .IN4(n456), .IN5(
          n483), .Q(tmp_sboxw[20]));
   AO221X1 U615 (.IN1(new_block[1]), .IN2(n451), .IN3(new_block[33]), .IN4(n455), .IN5(
          n484), .Q(tmp_sboxw[1]));
   AO22X1 U616 (.IN1(new_block[97]), .IN2(n453), .IN3(new_block[65]), .IN4(n449), .Q(n484)
          );
   AO221X1 U617 (.IN1(new_block[19]), .IN2(n451), .IN3(new_block[51]), .IN4(n455), .IN5(
          n485), .Q(tmp_sboxw[19]));
   AO22X1 U618 (.IN1(new_block[115]), .IN2(n453), .IN3(new_block[83]), .IN4(n449), .Q(n485)
          );
   AO221X1 U619 (.IN1(new_block[18]), .IN2(n451), .IN3(new_block[50]), .IN4(n455), .IN5(
          n486), .Q(tmp_sboxw[18]));
   AO22X1 U620 (.IN1(new_block[114]), .IN2(n453), .IN3(new_block[82]), .IN4(n449), .Q(n486)
          );
   AO221X1 U621 (.IN1(new_block[17]), .IN2(n451), .IN3(new_block[49]), .IN4(n455), .IN5(
          n487), .Q(tmp_sboxw[17]));
   AO22X1 U622 (.IN1(new_block[113]), .IN2(n453), .IN3(new_block[81]), .IN4(n449), .Q(n487)
          );
   AO221X1 U623 (.IN1(new_block[16]), .IN2(n451), .IN3(new_block[48]), .IN4(n455), .IN5(
          n488), .Q(tmp_sboxw[16]));
   AO22X1 U624 (.IN1(new_block[112]), .IN2(n453), .IN3(new_block[80]), .IN4(n449), .Q(n488)
          );
   AO221X1 U625 (.IN1(new_block[15]), .IN2(n451), .IN3(new_block[47]), .IN4(n455), .IN5(
          n489), .Q(tmp_sboxw[15]));
   AO22X1 U626 (.IN1(new_block[111]), .IN2(n453), .IN3(new_block[79]), .IN4(n449), .Q(n489)
          );
   AO221X1 U627 (.IN1(new_block[14]), .IN2(n451), .IN3(new_block[46]), .IN4(n455), .IN5(
          n490), .Q(tmp_sboxw[14]));
   AO22X1 U628 (.IN1(new_block[110]), .IN2(n453), .IN3(new_block[78]), .IN4(n449), .Q(n490)
          );
   AO221X1 U629 (.IN1(new_block[13]), .IN2(n451), .IN3(new_block[45]), .IN4(n455), .IN5(
          n491), .Q(tmp_sboxw[13]));
   AO22X1 U630 (.IN1(new_block[109]), .IN2(n453), .IN3(new_block[77]), .IN4(n449), .Q(n491)
          );
   AO221X1 U631 (.IN1(new_block[12]), .IN2(n451), .IN3(new_block[44]), .IN4(n455), .IN5(
          n492), .Q(tmp_sboxw[12]));
   AO22X1 U632 (.IN1(new_block[108]), .IN2(n453), .IN3(new_block[76]), .IN4(n449), .Q(n492)
          );
   AO221X1 U633 (.IN1(new_block[11]), .IN2(n451), .IN3(new_block[43]), .IN4(n455), .IN5(
          n493), .Q(tmp_sboxw[11]));
   AO22X1 U634 (.IN1(new_block[107]), .IN2(n453), .IN3(new_block[75]), .IN4(n449), .Q(n493)
          );
   AO221X1 U635 (.IN1(new_block[10]), .IN2(n451), .IN3(new_block[42]), .IN4(n455), .IN5(
          n494), .Q(tmp_sboxw[10]));
   AO22X1 U636 (.IN1(new_block[106]), .IN2(n453), .IN3(new_block[74]), .IN4(n449), .Q(n494)
          );
   AO221X1 U637 (.IN1(new_block[0]), .IN2(n451), .IN3(new_block[32]), .IN4(n455), .IN5(
          n495), .Q(tmp_sboxw[0]));
   AO22X1 U638 (.IN1(new_block[96]), .IN2(n453), .IN3(new_block[64]), .IN4(n449), .Q(n495)
          );
   AO221X1 U639 (.IN1(new_sboxw[31]), .IN2(n1081), .IN3(n409), .IN4(new_block[127]), .IN5(
          n501), .Q(n2006));
   OAI222X1 U640 (.IN1(n502), .IN2(n1231), .IN3(round_key[127]), .IN4(n503), .IN5(n504), .
          IN6(n1033), .QN(n501));
   XOR3X1 U642 (.IN1(n508), .IN2(n509), .IN3(n510), .Q(n507));
   XOR2X1 U643 (.IN1(n511), .IN2(n512), .Q(n510));
   XOR3X1 U645 (.IN1(n516), .IN2(n517), .IN3(n518), .Q(n515));
   AOI22X1 U646 (.IN1(n631), .IN2(block[127]), .IN3(new_block[127]), .IN4(n786), .QN(n503)
          );
   OA22X1 U647 (.IN1(new_block[127]), .IN2(n448), .IN3(block[127]), .IN4(n753), .Q(n502)
          );
   AO221X1 U648 (.IN1(new_sboxw[30]), .IN2(n1081), .IN3(n409), .IN4(new_block[126]), .IN5(
          n521), .Q(n2007));
   OAI222X1 U649 (.IN1(n522), .IN2(n1248), .IN3(round_key[126]), .IN4(n523), .IN5(n524), .
          IN6(n1033), .QN(n521));
   XOR3X1 U651 (.IN1(n527), .IN2(n1440), .IN3(n528), .Q(n526));
   XOR3X1 U653 (.IN1(n1537), .IN2(n531), .IN3(n532), .Q(n530));
   AOI22X1 U654 (.IN1(n646), .IN2(block[126]), .IN3(new_block[126]), .IN4(n832), .QN(n523)
          );
   OA22X1 U655 (.IN1(new_block[126]), .IN2(n448), .IN3(block[126]), .IN4(n753), .Q(n522)
          );
   AO221X1 U656 (.IN1(new_sboxw[29]), .IN2(n1081), .IN3(n409), .IN4(new_block[125]), .IN5(
          n533), .Q(n2008));
   OAI222X1 U657 (.IN1(n534), .IN2(n1262), .IN3(round_key[125]), .IN4(n535), .IN5(n536), .
          IN6(n1033), .QN(n533));
   XOR2X1 U660 (.IN1(n514), .IN2(n542), .Q(n541));
   XOR3X1 U661 (.IN1(n543), .IN2(n544), .IN3(n545), .Q(n537));
   XOR3X1 U662 (.IN1(n546), .IN2(n547), .IN3(n548), .Q(n545));
   AOI22X1 U663 (.IN1(n664), .IN2(block[125]), .IN3(new_block[125]), .IN4(n834), .QN(n535)
          );
   OA22X1 U664 (.IN1(new_block[125]), .IN2(n881), .IN3(block[125]), .IN4(n768), .Q(n534)
          );
   AO221X1 U665 (.IN1(new_sboxw[28]), .IN2(n1081), .IN3(n409), .IN4(new_block[124]), .IN5(
          n549), .Q(n2009));
   OAI222X1 U666 (.IN1(n550), .IN2(n1263), .IN3(round_key[124]), .IN4(n551), .IN5(n552), .
          IN6(n1033), .QN(n549));
   XOR3X1 U668 (.IN1(n555), .IN2(n514), .IN3(n556), .Q(n554));
   XOR2X1 U669 (.IN1(n557), .IN2(n532), .Q(n556));
   XNOR3X1 U671 (.IN1(n561), .IN2(n517), .IN3(n562), .Q(n560));
   AOI22X1 U672 (.IN1(n664), .IN2(block[124]), .IN3(new_block[124]), .IN4(n832), .QN(n551)
          );
   OA22X1 U673 (.IN1(new_block[124]), .IN2(n881), .IN3(block[124]), .IN4(n753), .Q(n550)
          );
   AO221X1 U674 (.IN1(new_sboxw[27]), .IN2(n1081), .IN3(n409), .IN4(new_block[123]), .IN5(
          n563), .Q(n2010));
   OAI222X1 U675 (.IN1(n564), .IN2(n1274), .IN3(round_key[123]), .IN4(n565), .IN5(n566), .
          IN6(n1033), .QN(n563));
   XOR3X1 U677 (.IN1(n569), .IN2(n570), .IN3(n571), .Q(n568));
   XOR2X1 U678 (.IN1(n572), .IN2(n573), .Q(n571));
   XOR3X1 U680 (.IN1(n577), .IN2(n578), .IN3(n579), .Q(n576));
   AOI22X1 U681 (.IN1(n679), .IN2(block[123]), .IN3(new_block[123]), .IN4(n834), .QN(n565)
          );
   OA22X1 U682 (.IN1(new_block[123]), .IN2(n519), .IN3(block[123]), .IN4(n768), .Q(n564)
          );
   AO221X1 U683 (.IN1(new_sboxw[26]), .IN2(n1081), .IN3(n409), .IN4(new_block[122]), .IN5(
          n580), .Q(n2011));
   OAI222X1 U684 (.IN1(n581), .IN2(n1275), .IN3(round_key[122]), .IN4(n582), .IN5(n583), .
          IN6(n1033), .QN(n580));
   XOR3X1 U686 (.IN1(n586), .IN2(n587), .IN3(n588), .Q(n585));
   XNOR3X1 U688 (.IN1(n592), .IN2(n593), .IN3(n594), .Q(n591));
   AOI22X1 U689 (.IN1(n697), .IN2(block[122]), .IN3(new_block[122]), .IN4(n435), .QN(n582)
          );
   OA22X1 U690 (.IN1(new_block[122]), .IN2(n850), .IN3(block[122]), .IN4(n753), .Q(n581)
          );
   AO221X1 U691 (.IN1(new_sboxw[25]), .IN2(n1081), .IN3(n409), .IN4(new_block[121]), .IN5(
          n595), .Q(n2012));
   OAI222X1 U692 (.IN1(n596), .IN2(n1276), .IN3(round_key[121]), .IN4(n597), .IN5(n598), .
          IN6(n1033), .QN(n595));
   XOR3X1 U694 (.IN1(n601), .IN2(n602), .IN3(n603), .Q(n600));
   XNOR2X1 U695 (.IN1(n604), .IN2(n605), .Q(n603));
   XOR3X1 U697 (.IN1(n609), .IN2(n610), .IN3(n611), .Q(n608));
   AOI22X1 U698 (.IN1(n679), .IN2(block[121]), .IN3(new_block[121]), .IN4(n437), .QN(n597)
          );
   OA22X1 U699 (.IN1(new_block[121]), .IN2(n897), .IN3(block[121]), .IN4(n753), .Q(n596)
          );
   AO221X1 U700 (.IN1(new_sboxw[24]), .IN2(n1081), .IN3(n409), .IN4(new_block[120]), .IN5(
          n612), .Q(n2013));
   OAI222X1 U701 (.IN1(n613), .IN2(n1286), .IN3(round_key[120]), .IN4(n614), .IN5(n615), .
          IN6(n1033), .QN(n612));
   XOR2X1 U702 (.IN1(n616), .IN2(n617), .Q(n615));
   XOR3X1 U705 (.IN1(n621), .IN2(n622), .IN3(n623), .Q(n616));
   XOR3X1 U706 (.IN1(n547), .IN2(n624), .IN3(n1416), .Q(n623));
   AOI22X1 U707 (.IN1(n679), .IN2(block[120]), .IN3(new_block[120]), .IN4(n434), .QN(n614)
          );
   OA22X1 U708 (.IN1(new_block[120]), .IN2(n850), .IN3(block[120]), .IN4(n753), .Q(n613)
          );
   AO221X1 U709 (.IN1(new_sboxw[23]), .IN2(n1081), .IN3(n679), .IN4(n626), .IN5(n627), .Q(
          n2014));
   OAI222X1 U710 (.IN1(n628), .IN2(n296), .IN3(n1287), .IN4(n629), .IN5(n630), .IN6(n1033)
          , .QN(n627));
   XOR3X1 U712 (.IN1(n633), .IN2(n634), .IN3(n635), .Q(n632));
   XOR3X1 U714 (.IN1(n638), .IN2(n639), .IN3(n640), .Q(n637));
   XOR2X1 U715 (.IN1(round_key[23]), .IN2(block[23]), .Q(n626));
   AO221X1 U716 (.IN1(new_sboxw[22]), .IN2(n1081), .IN3(n727), .IN4(n641), .IN5(n642), .Q(
          n2015));
   OAI222X1 U717 (.IN1(n643), .IN2(n298), .IN3(n1297), .IN4(n644), .IN5(n645), .IN6(n1022)
          , .QN(n642));
   XOR3X1 U719 (.IN1(n648), .IN2(n649), .IN3(n650), .Q(n647));
   XOR2X1 U720 (.IN1(n651), .IN2(n2200), .Q(n650));
   XOR3X1 U722 (.IN1(n655), .IN2(n656), .IN3(n657), .Q(n654));
   XOR2X1 U723 (.IN1(round_key[22]), .IN2(block[22]), .Q(n641));
   AO221X1 U724 (.IN1(new_sboxw[21]), .IN2(n1081), .IN3(n706), .IN4(n658), .IN5(n659), .Q(
          n2016));
   OAI222X1 U725 (.IN1(n660), .IN2(n300), .IN3(n1324), .IN4(n661), .IN5(n662), .IN6(n1022)
          , .QN(n659));
   XOR2X1 U728 (.IN1(n633), .IN2(n667), .Q(n665));
   XOR3X1 U729 (.IN1(n668), .IN2(n669), .IN3(n670), .Q(n663));
   XOR3X1 U730 (.IN1(n671), .IN2(n2181), .IN3(n672), .Q(n670));
   XOR2X1 U731 (.IN1(round_key[21]), .IN2(block[21]), .Q(n658));
   AO221X1 U732 (.IN1(new_sboxw[20]), .IN2(n1081), .IN3(n736), .IN4(n673), .IN5(n674), .Q(
          n2017));
   OAI222X1 U733 (.IN1(n675), .IN2(n302), .IN3(n1360), .IN4(n676), .IN5(n677), .IN6(n1022)
          , .QN(n674));
   XOR3X1 U735 (.IN1(n681), .IN2(n2219), .IN3(n682), .Q(n680));
   XOR2X1 U737 (.IN1(n2200), .IN2(n684), .Q(n683));
   XOR2X1 U738 (.IN1(round_key[20]), .IN2(block[20]), .Q(n673));
   AO221X1 U739 (.IN1(new_sboxw[19]), .IN2(n1087), .IN3(n736), .IN4(n685), .IN5(n686), .Q(
          n2018));
   OAI222X1 U740 (.IN1(n687), .IN2(n303), .IN3(n1371), .IN4(n688), .IN5(n689), .IN6(n1022)
          , .QN(n686));
   XOR3X1 U741 (.IN1(n690), .IN2(n691), .IN3(n692), .Q(n689));
   XOR3X1 U742 (.IN1(n693), .IN2(n2221), .IN3(n694), .Q(n692));
   XOR2X1 U745 (.IN1(round_key[19]), .IN2(block[19]), .Q(n685));
   AO221X1 U746 (.IN1(new_sboxw[18]), .IN2(n1087), .IN3(n706), .IN4(n699), .IN5(n700), .Q(
          n2019));
   OAI222X1 U747 (.IN1(n701), .IN2(n304), .IN3(n1372), .IN4(n702), .IN5(n703), .IN6(n1022)
          , .QN(n700));
   XOR3X1 U750 (.IN1(n710), .IN2(n711), .IN3(n712), .Q(n705));
   XOR2X1 U751 (.IN1(n713), .IN2(n714), .Q(n712));
   XOR2X1 U752 (.IN1(round_key[18]), .IN2(block[18]), .Q(n699));
   AO221X1 U753 (.IN1(new_sboxw[17]), .IN2(n1087), .IN3(n631), .IN4(n715), .IN5(n716), .Q(
          n2020));
   OAI222X1 U754 (.IN1(n717), .IN2(n305), .IN3(n1377), .IN4(n718), .IN5(n719), .IN6(n1022)
          , .QN(n716));
   XOR3X1 U755 (.IN1(n720), .IN2(n721), .IN3(n722), .Q(n719));
   XOR3X1 U756 (.IN1(n723), .IN2(n724), .IN3(n725), .Q(n722));
   XOR2X1 U759 (.IN1(round_key[17]), .IN2(block[17]), .Q(n715));
   AO221X1 U760 (.IN1(new_sboxw[16]), .IN2(n1087), .IN3(n727), .IN4(n729), .IN5(n730), .Q(
          n2021));
   OAI222X1 U761 (.IN1(n731), .IN2(n306), .IN3(n1382), .IN4(n732), .IN5(n733), .IN6(n1022)
          , .QN(n730));
   XOR3X1 U764 (.IN1(n740), .IN2(n2181), .IN3(n741), .Q(n735));
   XOR2X1 U765 (.IN1(n742), .IN2(n651), .Q(n741));
   XOR2X1 U766 (.IN1(n743), .IN2(n744), .Q(n734));
   XOR2X1 U767 (.IN1(round_key[16]), .IN2(block[16]), .Q(n729));
   AO221X1 U768 (.IN1(new_sboxw[15]), .IN2(n1087), .IN3(n727), .IN4(n745), .IN5(n746), .Q(
          n2022));
   OAI222X1 U769 (.IN1(n747), .IN2(n307), .IN3(n1390), .IN4(n748), .IN5(n749), .IN6(n1022)
          , .QN(n746));
   XOR3X1 U770 (.IN1(n750), .IN2(n751), .IN3(n752), .Q(n749));
   XOR3X1 U772 (.IN1(n755), .IN2(n756), .IN3(n757), .Q(n754));
   XOR2X1 U773 (.IN1(n758), .IN2(n759), .Q(n757));
   XOR2X1 U775 (.IN1(round_key[47]), .IN2(block[47]), .Q(n745));
   AO221X1 U776 (.IN1(new_sboxw[14]), .IN2(n1087), .IN3(n646), .IN4(n762), .IN5(n763), .Q(
          n2023));
   OAI222X1 U777 (.IN1(n764), .IN2(n313), .IN3(n1407), .IN4(n765), .IN5(n766), .IN6(n1022)
          , .QN(n763));
   XOR3X1 U780 (.IN1(n771), .IN2(n772), .IN3(n773), .Q(n770));
   XOR2X1 U781 (.IN1(n774), .IN2(n775), .Q(n773));
   XOR3X1 U782 (.IN1(n776), .IN2(n777), .IN3(n778), .Q(n769));
   XOR2X1 U783 (.IN1(round_key[46]), .IN2(block[46]), .Q(n762));
   AO221X1 U784 (.IN1(new_sboxw[13]), .IN2(n1087), .IN3(n706), .IN4(n779), .IN5(n780), .Q(
          n2024));
   OAI222X1 U785 (.IN1(n781), .IN2(n315), .IN3(n1450), .IN4(n782), .IN5(n783), .IN6(n1022)
          , .QN(n780));
   XOR3X1 U786 (.IN1(n755), .IN2(n767), .IN3(n784), .Q(n783));
   XOR2X1 U789 (.IN1(n790), .IN2(n1926), .Q(n787));
   XOR2X1 U791 (.IN1(round_key[45]), .IN2(block[45]), .Q(n779));
   AO221X1 U792 (.IN1(new_sboxw[12]), .IN2(n1087), .IN3(n697), .IN4(n794), .IN5(n795), .Q(
          n2025));
   OAI222X1 U793 (.IN1(n796), .IN2(n317), .IN3(n1460), .IN4(n797), .IN5(n798), .IN6(n1022)
          , .QN(n795));
   XNOR3X1 U795 (.IN1(n802), .IN2(n803), .IN3(n804), .Q(n801));
   XNOR3X1 U797 (.IN1(n805), .IN2(n806), .IN3(n807), .Q(n799));
   XOR2X1 U798 (.IN1(n808), .IN2(n809), .Q(n805));
   XOR2X1 U799 (.IN1(round_key[44]), .IN2(block[44]), .Q(n794));
   AO221X1 U800 (.IN1(new_sboxw[11]), .IN2(n1087), .IN3(n646), .IN4(n810), .IN5(n811), .Q(
          n2026));
   OAI222X1 U801 (.IN1(n812), .IN2(n318), .IN3(n1470), .IN4(n813), .IN5(n814), .IN6(n1022)
          , .QN(n811));
   XOR3X1 U803 (.IN1(n818), .IN2(n819), .IN3(n820), .Q(n817));
   XOR3X1 U805 (.IN1(n823), .IN2(n2156), .IN3(n824), .Q(n815));
   XOR2X1 U806 (.IN1(n825), .IN2(n826), .Q(n823));
   XOR2X1 U807 (.IN1(round_key[43]), .IN2(block[43]), .Q(n810));
   AO221X1 U808 (.IN1(new_sboxw[10]), .IN2(n1087), .IN3(n679), .IN4(n827), .IN5(n828), .Q(
          n2027));
   OAI222X1 U809 (.IN1(n829), .IN2(n319), .IN3(n1477), .IN4(n830), .IN5(n831), .IN6(n1022)
          , .QN(n828));
   XOR2X1 U814 (.IN1(n843), .IN2(n844), .Q(n842));
   XOR2X1 U815 (.IN1(round_key[42]), .IN2(block[42]), .Q(n827));
   AO221X1 U816 (.IN1(new_sboxw[9]), .IN2(n1087), .IN3(n664), .IN4(n845), .IN5(n846), .Q(
          n2028));
   OAI222X1 U817 (.IN1(n847), .IN2(n321), .IN3(n1486), .IN4(n848), .IN5(n849), .IN6(n1022)
          , .QN(n846));
   XNOR3X1 U819 (.IN1(n853), .IN2(n854), .IN3(n855), .Q(n852));
   XNOR2X1 U820 (.IN1(n839), .IN2(n856), .Q(n851));
   XOR2X1 U822 (.IN1(n860), .IN2(n861), .Q(n859));
   XOR2X1 U823 (.IN1(round_key[41]), .IN2(block[41]), .Q(n845));
   AO221X1 U824 (.IN1(new_sboxw[8]), .IN2(n1087), .IN3(n664), .IN4(n862), .IN5(n863), .Q(
          n2029));
   OAI222X1 U825 (.IN1(n864), .IN2(n322), .IN3(n1520), .IN4(n865), .IN5(n866), .IN6(n1022)
          , .QN(n863));
   XOR3X1 U827 (.IN1(n870), .IN2(n871), .IN3(n2158), .Q(n869));
   XOR3X1 U829 (.IN1(n872), .IN2(n873), .IN3(n874), .Q(n867));
   XOR2X1 U830 (.IN1(n875), .IN2(n791), .Q(n874));
   XOR2X1 U831 (.IN1(round_key[40]), .IN2(block[40]), .Q(n862));
   AO221X1 U832 (.IN1(new_sboxw[7]), .IN2(n1088), .IN3(n706), .IN4(n876), .IN5(n877), .Q(
          n2030));
   OAI222X1 U833 (.IN1(n878), .IN2(n323), .IN3(n1528), .IN4(n879), .IN5(n880), .IN6(n1008)
          , .QN(n877));
   XOR3X1 U835 (.IN1(n883), .IN2(n884), .IN3(n885), .Q(n882));
   XOR2X1 U836 (.IN1(n886), .IN2(n887), .Q(n885));
   XOR3X1 U838 (.IN1(n890), .IN2(n1614), .IN3(n891), .Q(n889));
   XOR2X1 U839 (.IN1(round_key[71]), .IN2(block[71]), .Q(n876));
   AO221X1 U840 (.IN1(new_sboxw[6]), .IN2(n1088), .IN3(n697), .IN4(n892), .IN5(n893), .Q(
          n2031));
   OAI222X1 U841 (.IN1(n894), .IN2(n326), .IN3(n1530), .IN4(n895), .IN5(n896), .IN6(n1008)
          , .QN(n893));
   XOR3X1 U843 (.IN1(n1614), .IN2(n899), .IN3(n900), .Q(n898));
   XOR2X1 U844 (.IN1(n1764), .IN2(n901), .Q(n900));
   XOR3X1 U846 (.IN1(n905), .IN2(n1623), .IN3(n906), .Q(n904));
   XOR2X1 U847 (.IN1(round_key[70]), .IN2(block[70]), .Q(n892));
   AO221X1 U848 (.IN1(new_sboxw[5]), .IN2(n1088), .IN3(n785), .IN4(n907), .IN5(n908), .Q(
          n2032));
   OAI222X1 U849 (.IN1(n909), .IN2(n328), .IN3(n1538), .IN4(n910), .IN5(n911), .IN6(n1008)
          , .QN(n908));
   XOR3X1 U852 (.IN1(n917), .IN2(n1634), .IN3(n918), .Q(n913));
   XOR2X1 U853 (.IN1(round_key[69]), .IN2(block[69]), .Q(n907));
   AO221X1 U854 (.IN1(new_sboxw[4]), .IN2(n1088), .IN3(n727), .IN4(n919), .IN5(n920), .Q(
          n2033));
   OAI222X1 U855 (.IN1(n921), .IN2(n330), .IN3(n1548), .IN4(n922), .IN5(n923), .IN6(n1008)
          , .QN(n920));
   XOR3X1 U858 (.IN1(n884), .IN2(n930), .IN3(n931), .Q(n925));
   XOR2X1 U859 (.IN1(n1634), .IN2(n1613), .Q(n931));
   XOR2X1 U860 (.IN1(round_key[68]), .IN2(block[68]), .Q(n919));
   AO221X1 U861 (.IN1(new_sboxw[3]), .IN2(n1088), .IN3(n785), .IN4(n932), .IN5(n933), .Q(
          n2034));
   OAI222X1 U862 (.IN1(n934), .IN2(n332), .IN3(n1556), .IN4(n935), .IN5(n936), .IN6(n1008)
          , .QN(n933));
   XOR3X1 U865 (.IN1(n943), .IN2(n944), .IN3(n945), .Q(n938));
   XOR2X1 U866 (.IN1(n946), .IN2(n947), .Q(n945));
   XOR2X1 U867 (.IN1(round_key[67]), .IN2(block[67]), .Q(n932));
   AO221X1 U868 (.IN1(new_sboxw[2]), .IN2(n1088), .IN3(n679), .IN4(n948), .IN5(n949), .Q(
          n2035));
   OAI222X1 U869 (.IN1(n950), .IN2(n333), .IN3(n1579), .IN4(n951), .IN5(n952), .IN6(n1008)
          , .QN(n949));
   XOR3X1 U870 (.IN1(n953), .IN2(n954), .IN3(n955), .Q(n952));
   XOR3X1 U871 (.IN1(n956), .IN2(n957), .IN3(n958), .Q(n955));
   XOR3X1 U872 (.IN1(n959), .IN2(n960), .IN3(n961), .Q(n954));
   XOR2X1 U873 (.IN1(n962), .IN2(n963), .Q(n961));
   XOR2X1 U874 (.IN1(round_key[66]), .IN2(block[66]), .Q(n948));
   AO221X1 U875 (.IN1(new_sboxw[1]), .IN2(n1088), .IN3(n785), .IN4(n964), .IN5(n965), .Q(
          n2036));
   OAI222X1 U876 (.IN1(n966), .IN2(n334), .IN3(n1594), .IN4(n967), .IN5(n968), .IN6(n1008)
          , .QN(n965));
   XOR3X1 U879 (.IN1(n963), .IN2(n975), .IN3(n976), .Q(n970));
   XNOR2X1 U880 (.IN1(n977), .IN2(n978), .Q(n976));
   XOR2X1 U881 (.IN1(round_key[65]), .IN2(block[65]), .Q(n964));
   AO221X1 U882 (.IN1(n567), .IN2(new_sboxw[31]), .IN3(n1), .IN4(new_block[95]), .IN5(n980)
          , .Q(n2037));
   OAI222X1 U883 (.IN1(n981), .IN2(n1606), .IN3(round_key[95]), .IN4(n982), .IN5(n983), .
          IN6(n1008), .QN(n980));
   XOR2X1 U886 (.IN1(n883), .IN2(n886), .Q(n986));
   XOR3X1 U887 (.IN1(n901), .IN2(n987), .IN3(n988), .Q(n984));
   XOR3X1 U888 (.IN1(n989), .IN2(n990), .IN3(n991), .Q(n988));
   AOI22X1 U889 (.IN1(n736), .IN2(block[95]), .IN3(new_block[95]), .IN4(n437), .QN(n982)
          );
   OA22X1 U890 (.IN1(new_block[95]), .IN2(n868), .IN3(block[95]), .IN4(n753), .Q(n981));
   AO221X1 U891 (.IN1(n567), .IN2(new_sboxw[30]), .IN3(n1), .IN4(new_block[94]), .IN5(n992)
          , .Q(n2038));
   OAI222X1 U892 (.IN1(n993), .IN2(n1615), .IN3(round_key[94]), .IN4(n994), .IN5(n995), .
          IN6(n1008), .QN(n992));
   XOR3X1 U894 (.IN1(n917), .IN2(n899), .IN3(n998), .Q(n997));
   XOR2X1 U895 (.IN1(n901), .IN2(n999), .Q(n998));
   XOR3X1 U897 (.IN1(n890), .IN2(n929), .IN3(n1003), .Q(n1002));
   AOI22X1 U898 (.IN1(n646), .IN2(block[94]), .IN3(new_block[94]), .IN4(n834), .QN(n994)
          );
   OA22X1 U899 (.IN1(new_block[94]), .IN2(n440), .IN3(block[94]), .IN4(n768), .Q(n993));
   AO221X1 U900 (.IN1(n567), .IN2(new_sboxw[29]), .IN3(n1), .IN4(new_block[93]), .IN5(
          n1004), .Q(n2039));
   OAI222X1 U901 (.IN1(n1005), .IN2(n1632), .IN3(round_key[93]), .IN4(n1006), .IN5(n1007)
          , .IN6(n1008), .QN(n1004));
   XOR3X1 U903 (.IN1(n917), .IN2(n930), .IN3(n1010), .Q(n1009));
   XOR2X1 U904 (.IN1(n1634), .IN2(n1011), .Q(n1010));
   XOR3X1 U906 (.IN1(n1015), .IN2(n1872), .IN3(n1016), .Q(n1014));
   AOI22X1 U907 (.IN1(n631), .IN2(block[93]), .IN3(new_block[93]), .IN4(n816), .QN(n1006)
          );
   OA22X1 U908 (.IN1(new_block[93]), .IN2(n447), .IN3(block[93]), .IN4(n768), .Q(n1005));
   AO221X1 U909 (.IN1(n567), .IN2(new_sboxw[28]), .IN3(n1), .IN4(new_block[92]), .IN5(
          n1017), .Q(n2040));
   OAI222X1 U910 (.IN1(n1018), .IN2(n1642), .IN3(round_key[92]), .IN4(n1019), .IN5(n1020)
          , .IN6(n1008), .QN(n1017));
   XOR2X1 U913 (.IN1(n1613), .IN2(n999), .Q(n1023));
   XOR3X1 U914 (.IN1(n1024), .IN2(n1025), .IN3(n1026), .Q(n1021));
   XOR3X1 U915 (.IN1(n1027), .IN2(n1892), .IN3(n1028), .Q(n1026));
   AOI22X1 U916 (.IN1(n631), .IN2(block[92]), .IN3(new_block[92]), .IN4(n816), .QN(n1019)
          );
   OA22X1 U917 (.IN1(new_block[92]), .IN2(n850), .IN3(block[92]), .IN4(n768), .Q(n1018));
   AO221X1 U918 (.IN1(n567), .IN2(new_sboxw[27]), .IN3(n1), .IN4(new_block[91]), .IN5(
          n1029), .Q(n2041));
   OAI222X1 U919 (.IN1(n1030), .IN2(n1651), .IN3(round_key[91]), .IN4(n1031), .IN5(n1032)
          , .IN6(n1008), .QN(n1029));
   XOR3X1 U921 (.IN1(n943), .IN2(n946), .IN3(n1035), .Q(n1034));
   XOR2X1 U922 (.IN1(n947), .IN2(n1036), .Q(n1035));
   XNOR3X1 U924 (.IN1(n1040), .IN2(n1041), .IN3(n1042), .Q(n1039));
   AOI22X1 U925 (.IN1(n646), .IN2(block[91]), .IN3(new_block[91]), .IN4(n786), .QN(n1031)
          );
   OA22X1 U926 (.IN1(new_block[91]), .IN2(n438), .IN3(block[91]), .IN4(n768), .Q(n1030));
   AO221X1 U927 (.IN1(n567), .IN2(new_sboxw[26]), .IN3(n1), .IN4(new_block[90]), .IN5(
          n1043), .Q(n2042));
   OAI222X1 U928 (.IN1(n1044), .IN2(n1661), .IN3(round_key[90]), .IN4(n1045), .IN5(n1046)
          , .IN6(n1008), .QN(n1043));
   XOR3X1 U930 (.IN1(n960), .IN2(n962), .IN3(n1049), .Q(n1048));
   XOR2X1 U931 (.IN1(n963), .IN2(n977), .Q(n1049));
   XOR3X1 U933 (.IN1(n1053), .IN2(n1054), .IN3(n1055), .Q(n1052));
   AOI22X1 U934 (.IN1(n646), .IN2(block[90]), .IN3(new_block[90]), .IN4(n435), .QN(n1045)
          );
   OA22X1 U935 (.IN1(new_block[90]), .IN2(n443), .IN3(block[90]), .IN4(n768), .Q(n1044));
   AO221X1 U936 (.IN1(n567), .IN2(new_sboxw[25]), .IN3(n1), .IN4(new_block[89]), .IN5(
          n1056), .Q(n2043));
   OAI222X1 U937 (.IN1(n1057), .IN2(n1674), .IN3(round_key[89]), .IN4(n1058), .IN5(n1059)
          , .IN6(n1008), .QN(n1056));
   XOR3X1 U939 (.IN1(n975), .IN2(n977), .IN3(n1062), .Q(n1061));
   XNOR2X1 U940 (.IN1(n978), .IN2(n1063), .Q(n1062));
   XOR3X1 U942 (.IN1(n956), .IN2(n1067), .IN3(n1068), .Q(n1066));
   AOI22X1 U943 (.IN1(n785), .IN2(block[89]), .IN3(new_block[89]), .IN4(n786), .QN(n1058)
          );
   OA22X1 U944 (.IN1(new_block[89]), .IN2(n442), .IN3(block[89]), .IN4(n768), .Q(n1057));
   AO221X1 U945 (.IN1(n567), .IN2(new_sboxw[24]), .IN3(n1), .IN4(new_block[88]), .IN5(
          n1069), .Q(n2044));
   OAI222X1 U946 (.IN1(n1070), .IN2(n1682), .IN3(round_key[88]), .IN4(n1071), .IN5(n1072)
          , .IN6(n1008), .QN(n1069));
   XOR2X1 U947 (.IN1(n1073), .IN2(n1074), .Q(n1072));
   XNOR3X1 U950 (.IN1(n1077), .IN2(n1078), .IN3(n1079), .Q(n1073));
   XOR3X1 U951 (.IN1(n905), .IN2(n1080), .IN3(n1771), .Q(n1079));
   AOI22X1 U952 (.IN1(n697), .IN2(block[88]), .IN3(new_block[88]), .IN4(n800), .QN(n1071)
          );
   OA22X1 U953 (.IN1(new_block[88]), .IN2(n868), .IN3(block[88]), .IN4(n753), .Q(n1070));
   AO221X1 U954 (.IN1(n567), .IN2(new_sboxw[23]), .IN3(n679), .IN4(n1082), .IN5(n1083), .Q(
          n2045));
   OAI222X1 U955 (.IN1(n1084), .IN2(n253), .IN3(n1691), .IN4(n1085), .IN5(n1086), .IN6(
          n996), .QN(n1083));
   XOR2X1 U960 (.IN1(round_key[119]), .IN2(block[119]), .Q(n1082));
   AO221X1 U961 (.IN1(n567), .IN2(new_sboxw[22]), .IN3(n697), .IN4(n1094), .IN5(n1095), .Q(
          n2046));
   OAI222X1 U962 (.IN1(n1096), .IN2(n256), .IN3(n1692), .IN4(n1097), .IN5(n1098), .IN6(
          n996), .QN(n1095));
   XOR3X1 U964 (.IN1(n1102), .IN2(n1537), .IN3(n1103), .Q(n1101));
   XOR2X1 U966 (.IN1(n1093), .IN2(n1399), .Q(n1104));
   XOR2X1 U968 (.IN1(round_key[118]), .IN2(block[118]), .Q(n1094));
   AO221X1 U969 (.IN1(n567), .IN2(new_sboxw[21]), .IN3(n631), .IN4(n1105), .IN5(n1106), .Q(
          n2047));
   OAI222X1 U970 (.IN1(n1107), .IN2(n258), .IN3(n1696), .IN4(n1108), .IN5(n1109), .IN6(
          n996), .QN(n1106));
   XOR3X1 U973 (.IN1(n1261), .IN2(n514), .IN3(n512), .Q(n1111));
   XOR2X1 U974 (.IN1(round_key[117]), .IN2(block[117]), .Q(n1105));
   AO221X1 U975 (.IN1(n567), .IN2(new_sboxw[20]), .IN3(n664), .IN4(n1115), .IN5(n1116), .Q(
          n2048));
   OAI222X1 U976 (.IN1(n1117), .IN2(n260), .IN3(n1709), .IN4(n1118), .IN5(n1119), .IN6(
          n996), .QN(n1116));
   XOR3X1 U977 (.IN1(n1120), .IN2(n1121), .IN3(n1122), .Q(n1119));
   XOR3X1 U978 (.IN1(n1123), .IN2(n1549), .IN3(n1124), .Q(n1122));
   XOR2X1 U981 (.IN1(round_key[116]), .IN2(block[116]), .Q(n1115));
   AO221X1 U982 (.IN1(n584), .IN2(new_sboxw[19]), .IN3(n646), .IN4(n1126), .IN5(n1127), .Q(
          n2049));
   OAI222X1 U983 (.IN1(n1128), .IN2(n261), .IN3(n1719), .IN4(n1129), .IN5(n1130), .IN6(
          n996), .QN(n1127));
   XOR3X1 U986 (.IN1(n569), .IN2(n1136), .IN3(n1137), .Q(n1132));
   XOR2X1 U987 (.IN1(n1392), .IN2(n573), .Q(n1137));
   XOR2X1 U988 (.IN1(round_key[115]), .IN2(block[115]), .Q(n1126));
   AO221X1 U989 (.IN1(n584), .IN2(new_sboxw[18]), .IN3(n631), .IN4(n1139), .IN5(n1140), .Q(
          n2050));
   OAI222X1 U990 (.IN1(n1141), .IN2(n262), .IN3(n1726), .IN4(n1142), .IN5(n1143), .IN6(
          n996), .QN(n1140));
   XOR3X1 U993 (.IN1(n1149), .IN2(n586), .IN3(n1150), .Q(n1145));
   XOR2X1 U994 (.IN1(n601), .IN2(n602), .Q(n1150));
   XOR2X1 U995 (.IN1(round_key[114]), .IN2(block[114]), .Q(n1139));
   AO221X1 U996 (.IN1(n584), .IN2(new_sboxw[17]), .IN3(n664), .IN4(n1151), .IN5(n1152), .Q(
          n2051));
   OAI222X1 U997 (.IN1(n1153), .IN2(n263), .IN3(n1738), .IN4(n1154), .IN5(n1155), .IN6(
          n996), .QN(n1152));
   XOR3X1 U998 (.IN1(n1156), .IN2(n1157), .IN3(n1158), .Q(n1155));
   XOR3X1 U999 (.IN1(n609), .IN2(n1159), .IN3(n1160), .Q(n1158));
   XOR3X1 U1000 (.IN1(n1161), .IN2(n601), .IN3(n1162), .Q(n1157));
   XOR2X1 U1001 (.IN1(n1391), .IN2(n605), .Q(n1162));
   XOR2X1 U1002 (.IN1(round_key[113]), .IN2(block[113]), .Q(n1151));
   AO221X1 U1003 (.IN1(n584), .IN2(new_sboxw[16]), .IN3(n664), .IN4(n1164), .IN5(n1165), .
          Q(n2052));
   OAI222X1 U1004 (.IN1(n1166), .IN2(n264), .IN3(n1744), .IN4(n1167), .IN5(n1168), .IN6(
          n996), .QN(n1165));
   XOR3X1 U1006 (.IN1(n624), .IN2(n610), .IN3(n611), .Q(n1171));
   XOR3X1 U1007 (.IN1(n508), .IN2(n1261), .IN3(n1172), .Q(n1170));
   XOR2X1 U1008 (.IN1(n511), .IN2(n539), .Q(n1172));
   XOR2X1 U1010 (.IN1(round_key[112]), .IN2(block[112]), .Q(n1164));
   AO221X1 U1011 (.IN1(n584), .IN2(new_sboxw[15]), .IN3(n706), .IN4(n1174), .IN5(n1175), .
          Q(n2053));
   OAI222X1 U1012 (.IN1(n1176), .IN2(n265), .IN3(n1752), .IN4(n1177), .IN5(n1178), .IN6(
          n996), .QN(n1175));
   XOR3X1 U1014 (.IN1(n655), .IN2(n1182), .IN3(n1183), .Q(n1181));
   XOR3X1 U1016 (.IN1(n639), .IN2(n740), .IN3(n1185), .Q(n1179));
   XOR2X1 U1017 (.IN1(n648), .IN2(n667), .Q(n1185));
   XOR2X1 U1018 (.IN1(round_key[15]), .IN2(block[15]), .Q(n1174));
   AO221X1 U1019 (.IN1(n584), .IN2(new_sboxw[14]), .IN3(n785), .IN4(n1186), .IN5(n1187), .
          Q(n2054));
   OAI222X1 U1020 (.IN1(n1188), .IN2(n270), .IN3(n1770), .IN4(n1189), .IN5(n1190), .IN6(
          n996), .QN(n1187));
   XOR3X1 U1024 (.IN1(n634), .IN2(n651), .IN3(n1197), .Q(n1191));
   XOR2X1 U1025 (.IN1(n684), .IN2(n656), .Q(n1197));
   XOR2X1 U1026 (.IN1(round_key[14]), .IN2(block[14]), .Q(n1186));
   AO221X1 U1027 (.IN1(n584), .IN2(new_sboxw[13]), .IN3(n706), .IN4(n1198), .IN5(n1199), .
          Q(n2055));
   OAI222X1 U1028 (.IN1(n1200), .IN2(n272), .IN3(n1779), .IN4(n1201), .IN5(n1202), .IN6(
          n996), .QN(n1199));
   XOR2X1 U1031 (.IN1(n671), .IN2(n1184), .Q(n1204));
   XOR2X1 U1034 (.IN1(round_key[13]), .IN2(block[13]), .Q(n1198));
   AO221X1 U1035 (.IN1(n584), .IN2(new_sboxw[12]), .IN3(n697), .IN4(n1211), .IN5(n1212), .
          Q(n2056));
   OAI222X1 U1036 (.IN1(n1213), .IN2(n274), .IN3(n1801), .IN4(n1214), .IN5(n1215), .IN6(
          n996), .QN(n1212));
   XOR2X1 U1041 (.IN1(n2183), .IN2(n667), .Q(n1222));
   XOR2X1 U1042 (.IN1(round_key[12]), .IN2(block[12]), .Q(n1211));
   AO221X1 U1043 (.IN1(n584), .IN2(new_sboxw[11]), .IN3(n697), .IN4(n1225), .IN5(n1226), .
          Q(n2057));
   OAI222X1 U1044 (.IN1(n1227), .IN2(n275), .IN3(n1817), .IN4(n1228), .IN5(n1229), .IN6(
          n996), .QN(n1226));
   XOR3X1 U1046 (.IN1(n1233), .IN2(n1234), .IN3(n1235), .Q(n1232));
   XOR3X1 U1048 (.IN1(n1238), .IN2(n1239), .IN3(n1240), .Q(n1230));
   XOR2X1 U1049 (.IN1(n696), .IN2(n1241), .Q(n1238));
   XOR2X1 U1050 (.IN1(round_key[11]), .IN2(block[11]), .Q(n1225));
   AO221X1 U1051 (.IN1(n584), .IN2(new_sboxw[10]), .IN3(n679), .IN4(n1242), .IN5(n1243), .
          Q(n2058));
   OAI222X1 U1052 (.IN1(n1244), .IN2(n276), .IN3(n1826), .IN4(n1245), .IN5(n1246), .IN6(
          n996), .QN(n1243));
   XOR3X1 U1054 (.IN1(n1250), .IN2(n1251), .IN3(n1252), .Q(n1249));
   XOR2X1 U1057 (.IN1(n713), .IN2(n1255), .Q(n1254));
   XOR2X1 U1058 (.IN1(round_key[10]), .IN2(block[10]), .Q(n1242));
   AO221X1 U1059 (.IN1(n584), .IN2(new_sboxw[9]), .IN3(n736), .IN4(n1256), .IN5(n1257), .Q(
          n2059));
   OAI222X1 U1060 (.IN1(n1258), .IN2(n277), .IN3(n1834), .IN4(n1259), .IN5(n1260), .IN6(
          n996), .QN(n1257));
   XOR2X1 U1065 (.IN1(n2198), .IN2(n739), .Q(n1267));
   XOR2X1 U1066 (.IN1(round_key[9]), .IN2(block[9]), .Q(n1256));
   AO221X1 U1067 (.IN1(n584), .IN2(new_sboxw[8]), .IN3(n697), .IN4(n1269), .IN5(n1270), .Q(
          n2060));
   OAI222X1 U1068 (.IN1(n1271), .IN2(n278), .IN3(n1842), .IN4(n1272), .IN5(n1273), .IN6(
          n985), .QN(n1270));
   XOR2X1 U1073 (.IN1(n742), .IN2(n649), .Q(n1280));
   XOR2X1 U1074 (.IN1(round_key[8]), .IN2(block[8]), .Q(n1269));
   AO221X1 U1075 (.IN1(n599), .IN2(new_sboxw[7]), .IN3(n736), .IN4(n1281), .IN5(n1282), .Q(
          n2061));
   OAI222X1 U1076 (.IN1(n1283), .IN2(n280), .IN3(n1852), .IN4(n1284), .IN5(n1285), .IN6(
          n985), .QN(n1282));
   XOR2X1 U1080 (.IN1(n756), .IN2(n790), .Q(n1291));
   XOR2X1 U1082 (.IN1(round_key[39]), .IN2(block[39]), .Q(n1281));
   AO221X1 U1083 (.IN1(n599), .IN2(new_sboxw[6]), .IN3(n679), .IN4(n1292), .IN5(n1293), .Q(
          n2062));
   OAI222X1 U1084 (.IN1(n1294), .IN2(n284), .IN3(n1862), .IN4(n1295), .IN5(n1296), .IN6(
          n985), .QN(n1293));
   XOR3X1 U1086 (.IN1(n1300), .IN2(n2171), .IN3(n1301), .Q(n1299));
   XOR3X1 U1087 (.IN1(n758), .IN2(n1926), .IN3(n1302), .Q(n1298));
   XOR2X1 U1088 (.IN1(n775), .IN2(n806), .Q(n1302));
   XOR2X1 U1090 (.IN1(round_key[38]), .IN2(block[38]), .Q(n1292));
   AO221X1 U1091 (.IN1(n599), .IN2(new_sboxw[5]), .IN3(n664), .IN4(n1304), .IN5(n1305), .Q(
          n2063));
   OAI222X1 U1092 (.IN1(n1306), .IN2(n286), .IN3(n1871), .IN4(n1307), .IN5(n1308), .IN6(
          n985), .QN(n1305));
   XOR3X1 U1094 (.IN1(n1312), .IN2(n2173), .IN3(n1313), .Q(n1311));
   XOR2X1 U1096 (.IN1(n1316), .IN2(n791), .Q(n1309));
   XOR2X1 U1097 (.IN1(round_key[37]), .IN2(block[37]), .Q(n1304));
   AO221X1 U1098 (.IN1(n599), .IN2(new_sboxw[4]), .IN3(n727), .IN4(n1317), .IN5(n1318), .Q(
          n2064));
   OAI222X1 U1099 (.IN1(n1319), .IN2(n288), .IN3(n1883), .IN4(n1320), .IN5(n1321), .IN6(
          n985), .QN(n1318));
   XOR3X1 U1102 (.IN1(n790), .IN2(n808), .IN3(n1327), .Q(n1323));
   XOR2X1 U1103 (.IN1(n809), .IN2(n1303), .Q(n1327));
   XOR2X1 U1104 (.IN1(round_key[36]), .IN2(block[36]), .Q(n1317));
   AO221X1 U1105 (.IN1(n599), .IN2(new_sboxw[3]), .IN3(n631), .IN4(n1328), .IN5(n1329), .Q(
          n2065));
   OAI222X1 U1106 (.IN1(n1330), .IN2(n289), .IN3(n1900), .IN4(n1331), .IN5(n1332), .IN6(
          n985), .QN(n1329));
   XOR3X1 U1107 (.IN1(n1333), .IN2(n1334), .IN3(n1335), .Q(n1332));
   XNOR3X1 U1108 (.IN1(n1336), .IN2(n822), .IN3(n1337), .Q(n1335));
   XOR3X1 U1109 (.IN1(n1338), .IN2(n825), .IN3(n1339), .Q(n1334));
   XOR2X1 U1110 (.IN1(n826), .IN2(n1340), .Q(n1339));
   XOR2X1 U1111 (.IN1(round_key[35]), .IN2(block[35]), .Q(n1328));
   AO221X1 U1112 (.IN1(n599), .IN2(new_sboxw[2]), .IN3(n646), .IN4(n1341), .IN5(n1342), .Q(
          n2066));
   OAI222X1 U1113 (.IN1(n1343), .IN2(n290), .IN3(n1901), .IN4(n1344), .IN5(n1345), .IN6(
          n985), .QN(n1342));
   XOR3X1 U1116 (.IN1(n1351), .IN2(n840), .IN3(n1352), .Q(n1347));
   XOR2X1 U1117 (.IN1(n841), .IN2(n857), .Q(n1352));
   XOR2X1 U1118 (.IN1(round_key[34]), .IN2(block[34]), .Q(n1341));
   AO221X1 U1119 (.IN1(n599), .IN2(new_sboxw[1]), .IN3(n727), .IN4(n1353), .IN5(n1354), .Q(
          n2067));
   OAI222X1 U1120 (.IN1(n1355), .IN2(n291), .IN3(n1902), .IN4(n1356), .IN5(n1357), .IN6(
          n985), .QN(n1354));
   XOR3X1 U1123 (.IN1(n857), .IN2(n843), .IN3(n1363), .Q(n1359));
   XNOR2X1 U1124 (.IN1(n858), .IN2(n1364), .Q(n1363));
   XOR2X1 U1125 (.IN1(round_key[33]), .IN2(block[33]), .Q(n1353));
   AO221X1 U1126 (.IN1(new_sboxw[0]), .IN2(n599), .IN3(n736), .IN4(n1365), .IN5(n1366), .Q(
          n2068));
   OAI222X1 U1127 (.IN1(n1367), .IN2(n292), .IN3(n1910), .IN4(n1368), .IN5(n1369), .IN6(
          n985), .QN(n1366));
   XOR2X1 U1131 (.IN1(n771), .IN2(n1926), .Q(n1314));
   XOR2X1 U1133 (.IN1(round_key[32]), .IN2(block[32]), .Q(n1365));
   AO221X1 U1135 (.IN1(n500), .IN2(new_sboxw[31]), .IN3(n463), .IN4(new_block[63]), .IN5(
          n1378), .Q(n2069));
   OAI222X1 U1136 (.IN1(n1379), .IN2(n1911), .IN3(round_key[63]), .IN4(n1380), .IN5(n1381)
          , .IN6(n985), .QN(n1378));
   XOR3X1 U1138 (.IN1(n775), .IN2(n875), .IN3(n1384), .Q(n1383));
   XOR3X1 U1139 (.IN1(n750), .IN2(n755), .IN3(n1912), .Q(n1384));
   XOR2X1 U1141 (.IN1(n2143), .IN2(n759), .Q(n1385));
   XOR2X1 U1142 (.IN1(n808), .IN2(n1926), .Q(n761));
   AOI22X1 U1143 (.IN1(n727), .IN2(block[63]), .IN3(new_block[63]), .IN4(n434), .QN(n1380)
          );
   OA22X1 U1144 (.IN1(new_block[63]), .IN2(n442), .IN3(block[63]), .IN4(n768), .Q(n1379)
          );
   AO221X1 U1145 (.IN1(n500), .IN2(new_sboxw[30]), .IN3(n463), .IN4(new_block[62]), .IN5(
          n1386), .Q(n2070));
   OAI222X1 U1146 (.IN1(n1387), .IN2(n1919), .IN3(round_key[62]), .IN4(n1388), .IN5(n1389)
          , .IN6(n985), .QN(n1386));
   XOR2X1 U1150 (.IN1(n758), .IN2(n1926), .Q(n1393));
   XOR2X1 U1153 (.IN1(n808), .IN2(n1303), .Q(n778));
   AOI22X1 U1154 (.IN1(n785), .IN2(block[62]), .IN3(new_block[62]), .IN4(n434), .QN(n1388)
          );
   OA22X1 U1155 (.IN1(new_block[62]), .IN2(n519), .IN3(block[62]), .IN4(n768), .Q(n1387)
          );
   AO221X1 U1156 (.IN1(n500), .IN2(new_sboxw[29]), .IN3(n463), .IN4(new_block[61]), .IN5(
          n1394), .Q(n2071));
   OAI222X1 U1157 (.IN1(n1395), .IN2(n1935), .IN3(round_key[61]), .IN4(n1396), .IN5(n1397)
          , .IN6(n985), .QN(n1394));
   XNOR2X1 U1160 (.IN1(n1315), .IN2(n806), .Q(n789));
   XOR2X1 U1161 (.IN1(n771), .IN2(n808), .Q(n1400));
   XOR3X1 U1162 (.IN1(n2147), .IN2(n793), .IN3(n1401), .Q(n1398));
   XOR3X1 U1163 (.IN1(n788), .IN2(n767), .IN3(n792), .Q(n1401));
   XNOR2X1 U1164 (.IN1(n1316), .IN2(n1303), .Q(n793));
   AOI22X1 U1165 (.IN1(n785), .IN2(block[61]), .IN3(new_block[61]), .IN4(n800), .QN(n1396)
          );
   OA22X1 U1166 (.IN1(new_block[61]), .IN2(n438), .IN3(block[61]), .IN4(n768), .Q(n1395)
          );
   AO221X1 U1167 (.IN1(n500), .IN2(new_sboxw[28]), .IN3(n463), .IN4(new_block[60]), .IN5(
          n1402), .Q(n2072));
   OAI222X1 U1168 (.IN1(n1403), .IN2(n1943), .IN3(round_key[60]), .IN4(n1404), .IN5(n1405)
          , .IN6(n985), .QN(n1402));
   XOR2X1 U1171 (.IN1(n1303), .IN2(n776), .Q(n1408));
   XOR3X1 U1172 (.IN1(n802), .IN2(n804), .IN3(n1409), .Q(n1406));
   XOR3X1 U1173 (.IN1(n807), .IN2(n755), .IN3(n803), .Q(n1409));
   XOR2X1 U1174 (.IN1(n1315), .IN2(n1410), .Q(n804));
   XOR2X1 U1175 (.IN1(n1316), .IN2(n1411), .Q(n802));
   AOI22X1 U1176 (.IN1(n736), .IN2(block[60]), .IN3(new_block[60]), .IN4(n800), .QN(n1404)
          );
   OA22X1 U1177 (.IN1(new_block[60]), .IN2(n446), .IN3(block[60]), .IN4(n768), .Q(n1403)
          );
   AO221X1 U1178 (.IN1(n500), .IN2(new_sboxw[27]), .IN3(n463), .IN4(new_block[59]), .IN5(
          n1412), .Q(n2073));
   OAI222X1 U1179 (.IN1(n1413), .IN2(n1953), .IN3(round_key[59]), .IN4(n1414), .IN5(n1415)
          , .IN6(n985), .QN(n1412));
   XOR3X1 U1181 (.IN1(n1338), .IN2(n826), .IN3(n1418), .Q(n1417));
   XOR2X1 U1182 (.IN1(n1340), .IN2(n1419), .Q(n1418));
   XOR3X1 U1184 (.IN1(n824), .IN2(n2175), .IN3(n820), .Q(n1420));
   XNOR2X1 U1185 (.IN1(n1421), .IN2(n1422), .Q(n819));
   XNOR2X1 U1186 (.IN1(n1423), .IN2(n1424), .Q(n818));
   AOI22X1 U1187 (.IN1(n697), .IN2(block[59]), .IN3(new_block[59]), .IN4(n832), .QN(n1414)
          );
   OA22X1 U1188 (.IN1(new_block[59]), .IN2(n436), .IN3(block[59]), .IN4(n768), .Q(n1413)
          );
   AO221X1 U1189 (.IN1(n500), .IN2(new_sboxw[26]), .IN3(n463), .IN4(new_block[58]), .IN5(
          n1425), .Q(n2074));
   OAI222X1 U1190 (.IN1(n1426), .IN2(n1962), .IN3(round_key[58]), .IN4(n1427), .IN5(n1428)
          , .IN6(n985), .QN(n1425));
   XOR2X1 U1191 (.IN1(n1429), .IN2(n1430), .Q(n1428));
   XOR3X1 U1192 (.IN1(n1351), .IN2(n841), .IN3(n1431), .Q(n1430));
   XOR2X1 U1193 (.IN1(n857), .IN2(n858), .Q(n1431));
   XOR3X1 U1194 (.IN1(n835), .IN2(n837), .IN3(n1432), .Q(n1429));
   XNOR3X1 U1195 (.IN1(n838), .IN2(n844), .IN3(n836), .Q(n1432));
   XNOR2X1 U1196 (.IN1(n2155), .IN2(n1433), .Q(n837));
   XNOR2X1 U1197 (.IN1(n1364), .IN2(n1434), .Q(n835));
   AOI22X1 U1198 (.IN1(n631), .IN2(block[58]), .IN3(new_block[58]), .IN4(n832), .QN(n1427)
          );
   OA22X1 U1199 (.IN1(new_block[58]), .IN2(n868), .IN3(block[58]), .IN4(n768), .Q(n1426)
          );
   AO221X1 U1200 (.IN1(n500), .IN2(new_sboxw[25]), .IN3(n463), .IN4(new_block[57]), .IN5(
          n1435), .Q(n2075));
   OAI222X1 U1201 (.IN1(n1436), .IN2(n1970), .IN3(round_key[57]), .IN4(n1437), .IN5(n1438)
          , .IN6(n979), .QN(n1435));
   XNOR2X1 U1204 (.IN1(n1364), .IN2(n1442), .Q(n1441));
   XOR3X1 U1205 (.IN1(n853), .IN2(n855), .IN3(n1443), .Q(n1439));
   XNOR3X1 U1206 (.IN1(n839), .IN2(n861), .IN3(n854), .Q(n1443));
   XNOR2X1 U1207 (.IN1(n2158), .IN2(n1433), .Q(n855));
   XOR2X1 U1208 (.IN1(n871), .IN2(n1434), .Q(n853));
   AOI22X1 U1209 (.IN1(n706), .IN2(block[57]), .IN3(new_block[57]), .IN4(n833), .QN(n1437)
          );
   OA22X1 U1210 (.IN1(new_block[57]), .IN2(n436), .IN3(block[57]), .IN4(n753), .Q(n1436)
          );
   AO221X1 U1211 (.IN1(n500), .IN2(new_sboxw[24]), .IN3(n463), .IN4(new_block[56]), .IN5(
          n1444), .Q(n2076));
   OAI222X1 U1212 (.IN1(n1445), .IN2(n1977), .IN3(round_key[56]), .IN4(n1446), .IN5(n1447)
          , .IN6(n979), .QN(n1444));
   XOR2X1 U1213 (.IN1(n1448), .IN2(n1449), .Q(n1447));
   XOR3X1 U1216 (.IN1(n870), .IN2(n871), .IN3(n1451), .Q(n1448));
   XOR3X1 U1217 (.IN1(n767), .IN2(n872), .IN3(n2158), .Q(n1451));
   AOI22X1 U1218 (.IN1(n727), .IN2(block[56]), .IN3(new_block[56]), .IN4(n914), .QN(n1446)
          );
   OA22X1 U1219 (.IN1(new_block[56]), .IN2(n519), .IN3(block[56]), .IN4(n768), .Q(n1445)
          );
   AO221X1 U1220 (.IN1(n500), .IN2(new_sboxw[23]), .IN3(n631), .IN4(n1454), .IN5(n1455), .
          Q(n2077));
   OAI222X1 U1221 (.IN1(n1456), .IN2(n209), .IN3(n1988), .IN4(n1457), .IN5(n1458), .IN6(
          n979), .QN(n1455));
   XOR2X1 U1224 (.IN1(n887), .IN2(n1634), .Q(n1461));
   XOR2X1 U1225 (.IN1(n930), .IN2(n917), .Q(n887));
   XOR3X1 U1226 (.IN1(n888), .IN2(n899), .IN3(n1462), .Q(n1459));
   XOR3X1 U1227 (.IN1(n990), .IN2(n901), .IN3(n891), .Q(n1462));
   XOR2X1 U1228 (.IN1(n1892), .IN2(n905), .Q(n891));
   XOR2X1 U1229 (.IN1(round_key[87]), .IN2(block[87]), .Q(n1454));
   AO221X1 U1230 (.IN1(n500), .IN2(new_sboxw[22]), .IN3(n631), .IN4(n1463), .IN5(n1464), .
          Q(n2078));
   OAI222X1 U1231 (.IN1(n1465), .IN2(n211), .IN3(n2144), .IN4(n1466), .IN5(n1467), .IN6(
          n979), .QN(n1464));
   XOR2X1 U1232 (.IN1(n1468), .IN2(n1469), .Q(n1467));
   XOR3X1 U1235 (.IN1(n902), .IN2(n903), .IN3(n1471), .Q(n1468));
   XOR3X1 U1236 (.IN1(n890), .IN2(n1011), .IN3(n906), .Q(n1471));
   XOR2X1 U1237 (.IN1(n1892), .IN2(n929), .Q(n906));
   XOR2X1 U1239 (.IN1(round_key[86]), .IN2(block[86]), .Q(n1463));
   AO221X1 U1240 (.IN1(n500), .IN2(new_sboxw[21]), .IN3(n646), .IN4(n1472), .IN5(n1473), .
          Q(n2079));
   OAI222X1 U1241 (.IN1(n1474), .IN2(n213), .IN3(n2146), .IN4(n1475), .IN5(n1476), .IN6(
          n979), .QN(n1473));
   XOR3X1 U1243 (.IN1(n915), .IN2(n1872), .IN3(n916), .Q(n1478));
   XOR2X1 U1244 (.IN1(n1013), .IN2(n999), .Q(n916));
   XOR2X1 U1245 (.IN1(n1015), .IN2(n929), .Q(n915));
   XOR2X1 U1248 (.IN1(round_key[85]), .IN2(block[85]), .Q(n1472));
   AO221X1 U1249 (.IN1(n500), .IN2(new_sboxw[20]), .IN3(n664), .IN4(n1481), .IN5(n1482), .
          Q(n2080));
   OAI222X1 U1250 (.IN1(n1483), .IN2(n215), .IN3(n2148), .IN4(n1484), .IN5(n1485), .IN6(
          n979), .QN(n1482));
   XOR3X1 U1252 (.IN1(n927), .IN2(n1892), .IN3(n928), .Q(n1487));
   XOR2X1 U1256 (.IN1(n1764), .IN2(n999), .Q(n1488));
   XOR2X1 U1257 (.IN1(n1489), .IN2(n1490), .Q(n924));
   XOR2X1 U1258 (.IN1(round_key[84]), .IN2(block[84]), .Q(n1481));
   AO221X1 U1259 (.IN1(n506), .IN2(new_sboxw[19]), .IN3(n785), .IN4(n1491), .IN5(n1492), .
          Q(n2081));
   OAI222X1 U1260 (.IN1(n1493), .IN2(n216), .IN3(n2150), .IN4(n1494), .IN5(n1495), .IN6(
          n979), .QN(n1492));
   XOR2X1 U1263 (.IN1(n1038), .IN2(n1498), .Q(n942));
   XOR2X1 U1264 (.IN1(n1040), .IN2(n1499), .Q(n940));
   XOR3X1 U1265 (.IN1(n943), .IN2(n944), .IN3(n1500), .Q(n1496));
   XOR2X1 U1266 (.IN1(n1760), .IN2(n1036), .Q(n1500));
   XOR2X1 U1267 (.IN1(n1502), .IN2(n1503), .Q(n937));
   XOR2X1 U1268 (.IN1(round_key[83]), .IN2(block[83]), .Q(n1491));
   AO221X1 U1269 (.IN1(n506), .IN2(new_sboxw[18]), .IN3(n706), .IN4(n1504), .IN5(n1505), .
          Q(n2082));
   OAI222X1 U1270 (.IN1(n1506), .IN2(n217), .IN3(n2151), .IN4(n1507), .IN5(n1508), .IN6(
          n979), .QN(n1505));
   XOR3X1 U1271 (.IN1(n953), .IN2(n1509), .IN3(n1510), .Q(n1508));
   XOR3X1 U1272 (.IN1(n1053), .IN2(n957), .IN3(n958), .Q(n1510));
   XNOR2X1 U1273 (.IN1(n1063), .IN2(n1050), .Q(n958));
   XOR2X1 U1274 (.IN1(n972), .IN2(n1054), .Q(n957));
   XOR3X1 U1275 (.IN1(n959), .IN2(n960), .IN3(n1511), .Q(n1509));
   XOR2X1 U1276 (.IN1(n975), .IN2(n977), .Q(n1511));
   XOR2X1 U1277 (.IN1(n1512), .IN2(n1513), .Q(n953));
   XOR2X1 U1278 (.IN1(round_key[82]), .IN2(block[82]), .Q(n1504));
   AO221X1 U1279 (.IN1(n506), .IN2(new_sboxw[17]), .IN3(n697), .IN4(n1514), .IN5(n1515), .
          Q(n2083));
   OAI222X1 U1280 (.IN1(n1516), .IN2(n218), .IN3(n2152), .IN4(n1517), .IN5(n1518), .IN6(
          n979), .QN(n1515));
   XOR2X1 U1283 (.IN1(n1863), .IN2(n1054), .Q(n974));
   XOR2X1 U1284 (.IN1(n1064), .IN2(n1050), .Q(n973));
   XOR3X1 U1285 (.IN1(n963), .IN2(n975), .IN3(n1521), .Q(n1519));
   XNOR2X1 U1286 (.IN1(n1522), .IN2(n1063), .Q(n1521));
   XOR2X1 U1287 (.IN1(n1078), .IN2(n1771), .Q(n969));
   XOR2X1 U1288 (.IN1(round_key[81]), .IN2(block[81]), .Q(n1514));
   AO221X1 U1289 (.IN1(n506), .IN2(new_sboxw[16]), .IN3(n697), .IN4(n1523), .IN5(n1524), .
          Q(n2084));
   OAI222X1 U1290 (.IN1(n1525), .IN2(n219), .IN3(n2153), .IN4(n1526), .IN5(n1527), .IN6(
          n979), .QN(n1524));
   XOR3X1 U1293 (.IN1(n883), .IN2(n886), .IN3(n918), .Q(n1529));
   XOR2X1 U1294 (.IN1(n1623), .IN2(n1011), .Q(n918));
   XOR2X1 U1296 (.IN1(round_key[80]), .IN2(block[80]), .Q(n1523));
   AO221X1 U1297 (.IN1(n506), .IN2(new_sboxw[15]), .IN3(n631), .IN4(n1532), .IN5(n1533), .
          Q(n2085));
   OAI222X1 U1298 (.IN1(n1534), .IN2(n222), .IN3(n2154), .IN4(n1535), .IN5(n1536), .IN6(
          n979), .QN(n1533));
   XOR2X1 U1301 (.IN1(n1288), .IN2(n512), .Q(n1540));
   XOR2X1 U1302 (.IN1(n539), .IN2(n555), .Q(n512));
   XOR2X1 U1303 (.IN1(n540), .IN2(n1261), .Q(n513));
   XOR2X1 U1306 (.IN1(round_key[111]), .IN2(block[111]), .Q(n1532));
   AO221X1 U1307 (.IN1(n506), .IN2(new_sboxw[14]), .IN3(n646), .IN4(n1542), .IN5(n1543), .
          Q(n2086));
   OAI222X1 U1308 (.IN1(n1544), .IN2(n225), .IN3(n2157), .IN4(n1545), .IN5(n1546), .IN6(
          n979), .QN(n1543));
   XOR3X1 U1309 (.IN1(n1541), .IN2(n531), .IN3(n1547), .Q(n1546));
   XOR2X1 U1313 (.IN1(n539), .IN2(n509), .Q(n1550));
   XNOR2X1 U1315 (.IN1(n540), .IN2(n557), .Q(n529));
   XOR2X1 U1316 (.IN1(round_key[110]), .IN2(block[110]), .Q(n1542));
   AO221X1 U1317 (.IN1(n506), .IN2(new_sboxw[13]), .IN3(n706), .IN4(n1551), .IN5(n1552), .
          Q(n2087));
   OAI222X1 U1318 (.IN1(n1553), .IN2(n227), .IN3(n2160), .IN4(n1554), .IN5(n1555), .IN6(
          n979), .QN(n1552));
   XOR3X1 U1321 (.IN1(n1559), .IN2(n1348), .IN3(n544), .Q(n1558));
   XNOR2X1 U1322 (.IN1(n1560), .IN2(n557), .Q(n544));
   XOR2X1 U1323 (.IN1(n555), .IN2(n1261), .Q(n1559));
   XNOR3X1 U1324 (.IN1(n548), .IN2(n546), .IN3(n543), .Q(n1557));
   XOR2X1 U1325 (.IN1(n1561), .IN2(n1562), .Q(n543));
   XOR2X1 U1326 (.IN1(round_key[109]), .IN2(block[109]), .Q(n1551));
   AO221X1 U1327 (.IN1(n506), .IN2(new_sboxw[12]), .IN3(n736), .IN4(n1563), .IN5(n1564), .
          Q(n2088));
   OAI222X1 U1328 (.IN1(n1565), .IN2(n229), .IN3(n2161), .IN4(n1566), .IN5(n1567), .IN6(
          n979), .QN(n1564));
   XOR3X1 U1331 (.IN1(n1571), .IN2(n1562), .IN3(n558), .Q(n1570));
   XNOR2X1 U1332 (.IN1(n1560), .IN2(n1572), .Q(n558));
   XOR2X1 U1333 (.IN1(n540), .IN2(n514), .Q(n1571));
   XNOR3X1 U1334 (.IN1(n562), .IN2(n561), .IN3(n559), .Q(n1569));
   XOR2X1 U1335 (.IN1(n1561), .IN2(n1573), .Q(n559));
   XOR2X1 U1336 (.IN1(round_key[108]), .IN2(block[108]), .Q(n1563));
   AO221X1 U1337 (.IN1(n506), .IN2(new_sboxw[11]), .IN3(n646), .IN4(n1574), .IN5(n1575), .
          Q(n2089));
   OAI222X1 U1338 (.IN1(n1576), .IN2(n230), .IN3(n2162), .IN4(n1577), .IN5(n1578), .IN6(
          n979), .QN(n1575));
   XOR3X1 U1341 (.IN1(n1582), .IN2(n1138), .IN3(n575), .Q(n1581));
   XNOR2X1 U1342 (.IN1(n1583), .IN2(n1584), .Q(n575));
   XOR2X1 U1343 (.IN1(n1136), .IN2(n570), .Q(n1582));
   XNOR3X1 U1344 (.IN1(n579), .IN2(n577), .IN3(n574), .Q(n1580));
   XNOR2X1 U1345 (.IN1(n1585), .IN2(n1586), .Q(n574));
   XOR2X1 U1346 (.IN1(round_key[107]), .IN2(block[107]), .Q(n1574));
   AO221X1 U1347 (.IN1(n506), .IN2(new_sboxw[10]), .IN3(n679), .IN4(n1588), .IN5(n1589), .
          Q(n2090));
   OAI222X1 U1348 (.IN1(n1590), .IN2(n231), .IN3(n2163), .IN4(n1591), .IN5(n1592), .IN6(
          n971), .QN(n1589));
   XOR3X1 U1349 (.IN1(n592), .IN2(n609), .IN3(n1593), .Q(n1592));
   XOR2X1 U1352 (.IN1(n604), .IN2(n1597), .Q(n589));
   XOR2X1 U1353 (.IN1(n1149), .IN2(n587), .Q(n1596));
   XNOR2X1 U1355 (.IN1(n1163), .IN2(n1598), .Q(n590));
   XOR2X1 U1356 (.IN1(round_key[106]), .IN2(block[106]), .Q(n1588));
   AO221X1 U1357 (.IN1(n506), .IN2(new_sboxw[9]), .IN3(n727), .IN4(n1599), .IN5(n1600), .Q(
          n2091));
   OAI222X1 U1358 (.IN1(n1601), .IN2(n232), .IN3(n2164), .IN4(n1602), .IN5(n1603), .IN6(
          n971), .QN(n1600));
   XNOR3X1 U1359 (.IN1(n609), .IN2(n1604), .IN3(n1605), .Q(n1603));
   XOR3X1 U1361 (.IN1(n588), .IN2(n1163), .IN3(n606), .Q(n1607));
   XNOR2X1 U1362 (.IN1(n622), .IN2(n1597), .Q(n606));
   XOR2X1 U1363 (.IN1(n1161), .IN2(n602), .Q(n588));
   XNOR2X1 U1365 (.IN1(n1416), .IN2(n1598), .Q(n607));
   XOR2X1 U1366 (.IN1(round_key[105]), .IN2(block[105]), .Q(n1599));
   AO221X1 U1367 (.IN1(n506), .IN2(new_sboxw[8]), .IN3(n697), .IN4(n1608), .IN5(n1609), .Q(
          n2092));
   OAI222X1 U1368 (.IN1(n1610), .IN2(n233), .IN3(n2165), .IN4(n1611), .IN5(n1612), .IN6(
          n971), .QN(n1609));
   XOR2X1 U1373 (.IN1(n511), .IN2(n542), .Q(n1617));
   XOR2X1 U1374 (.IN1(round_key[104]), .IN2(block[104]), .Q(n1608));
   AO221X1 U1375 (.IN1(n525), .IN2(new_sboxw[7]), .IN3(n697), .IN4(n1618), .IN5(n1619), .Q(
          n2093));
   OAI222X1 U1376 (.IN1(n1620), .IN2(n234), .IN3(n2166), .IN4(n1621), .IN5(n1622), .IN6(
          n971), .QN(n1619));
   XOR3X1 U1378 (.IN1(n742), .IN2(n633), .IN3(n1625), .Q(n1624));
   XOR2X1 U1379 (.IN1(n2183), .IN2(n636), .Q(n1625));
   XOR2X1 U1380 (.IN1(n667), .IN2(n649), .Q(n636));
   XOR3X1 U1382 (.IN1(n655), .IN2(n656), .IN3(n640), .Q(n1626));
   XOR2X1 U1383 (.IN1(n2219), .IN2(n671), .Q(n640));
   XOR2X1 U1384 (.IN1(round_key[7]), .IN2(block[7]), .Q(n1618));
   AO221X1 U1385 (.IN1(n525), .IN2(new_sboxw[6]), .IN3(n727), .IN4(n1627), .IN5(n1628), .Q(
          n2094));
   OAI222X1 U1386 (.IN1(n1629), .IN2(n237), .IN3(n2168), .IN4(n1630), .IN5(n1631), .IN6(
          n971), .QN(n1628));
   XOR2X1 U1389 (.IN1(n2219), .IN2(n2213), .Q(n657));
   XOR3X1 U1390 (.IN1(n648), .IN2(n634), .IN3(n1635), .Q(n1633));
   XOR2X1 U1391 (.IN1(n2200), .IN2(n653), .Q(n1635));
   XOR2X1 U1394 (.IN1(round_key[6]), .IN2(block[6]), .Q(n1627));
   AO221X1 U1395 (.IN1(n525), .IN2(new_sboxw[5]), .IN3(n736), .IN4(n1636), .IN5(n1637), .Q(
          n2095));
   OAI222X1 U1396 (.IN1(n1638), .IN2(n239), .IN3(n2170), .IN4(n1639), .IN5(n1640), .IN6(
          n971), .QN(n1637));
   XOR3X1 U1399 (.IN1(n668), .IN2(n669), .IN3(n1644), .Q(n1641));
   XOR3X1 U1400 (.IN1(n1184), .IN2(n2181), .IN3(n672), .Q(n1644));
   XOR2X1 U1401 (.IN1(n1207), .IN2(n2213), .Q(n672));
   XOR2X1 U1402 (.IN1(n1210), .IN2(n684), .Q(n668));
   XOR2X1 U1403 (.IN1(round_key[5]), .IN2(block[5]), .Q(n1636));
   AO221X1 U1404 (.IN1(n525), .IN2(new_sboxw[4]), .IN3(n706), .IN4(n1645), .IN5(n1646), .Q(
          n2096));
   OAI222X1 U1405 (.IN1(n1647), .IN2(n241), .IN3(n2172), .IN4(n1648), .IN5(n1649), .IN6(
          n971), .QN(n1646));
   XOR3X1 U1410 (.IN1(n633), .IN2(n2183), .IN3(n1652), .Q(n1650));
   XOR2X1 U1411 (.IN1(n667), .IN2(n653), .Q(n1652));
   XOR2X1 U1412 (.IN1(n1653), .IN2(n1654), .Q(n678));
   XOR2X1 U1413 (.IN1(round_key[4]), .IN2(block[4]), .Q(n1645));
   AO221X1 U1414 (.IN1(n525), .IN2(new_sboxw[3]), .IN3(n736), .IN4(n1655), .IN5(n1656), .Q(
          n2097));
   OAI222X1 U1415 (.IN1(n1657), .IN2(n243), .IN3(n2174), .IN4(n1658), .IN5(n1659), .IN6(
          n971), .QN(n1656));
   XOR2X1 U1418 (.IN1(n1240), .IN2(n1662), .Q(n694));
   XOR2X1 U1419 (.IN1(n1234), .IN2(n1663), .Q(n693));
   XOR3X1 U1420 (.IN1(n695), .IN2(n696), .IN3(n1664), .Q(n1660));
   XOR2X1 U1421 (.IN1(n1241), .IN2(n1665), .Q(n1664));
   XOR2X1 U1422 (.IN1(n1666), .IN2(n1667), .Q(n690));
   XOR2X1 U1423 (.IN1(round_key[3]), .IN2(block[3]), .Q(n1655));
   AO221X1 U1424 (.IN1(n525), .IN2(new_sboxw[2]), .IN3(n706), .IN4(n1668), .IN5(n1669), .Q(
          n2098));
   OAI222X1 U1425 (.IN1(n1670), .IN2(n244), .IN3(n2176), .IN4(n1671), .IN5(n1672), .IN6(
          n971), .QN(n1669));
   XNOR2X1 U1428 (.IN1(n728), .IN2(n1255), .Q(n709));
   XOR2X1 U1429 (.IN1(n1266), .IN2(n1250), .Q(n708));
   XOR3X1 U1430 (.IN1(n710), .IN2(n711), .IN3(n1675), .Q(n1673));
   XOR2X1 U1431 (.IN1(n1253), .IN2(n726), .Q(n1675));
   XOR2X1 U1432 (.IN1(n1676), .IN2(n635), .Q(n704));
   XOR2X1 U1433 (.IN1(round_key[2]), .IN2(block[2]), .Q(n1668));
   AO221X1 U1434 (.IN1(n525), .IN2(new_sboxw[1]), .IN3(n706), .IN4(n1677), .IN5(n1678), .Q(
          n2099));
   OAI222X1 U1435 (.IN1(n1679), .IN2(n245), .IN3(n2177), .IN4(n1680), .IN5(n1681), .IN6(
          n971), .QN(n1678));
   XOR3X1 U1437 (.IN1(n1266), .IN2(n724), .IN3(n725), .Q(n1683));
   XNOR2X1 U1438 (.IN1(n739), .IN2(n1255), .Q(n725));
   XOR2X1 U1439 (.IN1(n738), .IN2(n1250), .Q(n724));
   XNOR2X1 U1441 (.IN1(n714), .IN2(n1685), .Q(n1684));
   XOR2X1 U1442 (.IN1(n1277), .IN2(n2202), .Q(n720));
   XOR2X1 U1443 (.IN1(round_key[1]), .IN2(block[1]), .Q(n1677));
   AO221X1 U1444 (.IN1(n525), .IN2(new_sboxw[0]), .IN3(n727), .IN4(n1686), .IN5(n1687), .Q(
          n2100));
   OAI222X1 U1445 (.IN1(n1688), .IN2(n246), .IN3(n2178), .IN4(n1689), .IN5(n1690), .IN6(
          n971), .QN(n1687));
   XOR2X1 U1449 (.IN1(n639), .IN2(n651), .Q(n1694));
   XOR2X1 U1451 (.IN1(round_key[0]), .IN2(block[0]), .Q(n1686));
   AO221X1 U1453 (.IN1(n459), .IN2(new_sboxw[31]), .IN3(n144), .IN4(new_block[31]), .IN5(
          n1697), .Q(n2101));
   OAI222X1 U1454 (.IN1(n1698), .IN2(n2179), .IN3(round_key[31]), .IN4(n1699), .IN5(n1700)
          , .IN6(n971), .QN(n1697));
   XOR2X1 U1455 (.IN1(n1701), .IN2(n1702), .Q(n1700));
   XOR3X1 U1458 (.IN1(n656), .IN2(n1182), .IN3(n1704), .Q(n1701));
   XOR3X1 U1459 (.IN1(n638), .IN2(n1184), .IN3(n1183), .Q(n1704));
   XOR2X1 U1460 (.IN1(n2207), .IN2(n651), .Q(n1183));
   XOR2X1 U1461 (.IN1(n2183), .IN2(n2181), .Q(n1182));
   AOI22X1 U1462 (.IN1(n736), .IN2(block[31]), .IN3(new_block[31]), .IN4(n914), .QN(n1699)
          );
   OA22X1 U1463 (.IN1(new_block[31]), .IN2(n850), .IN3(block[31]), .IN4(n768), .Q(n1698)
          );
   AO221X1 U1464 (.IN1(n459), .IN2(new_sboxw[30]), .IN3(n144), .IN4(new_block[30]), .IN5(
          n1705), .Q(n2102));
   OAI222X1 U1465 (.IN1(n1706), .IN2(n2180), .IN3(round_key[30]), .IN4(n1707), .IN5(n1708)
          , .IN6(n971), .QN(n1705));
   XOR3X1 U1467 (.IN1(n648), .IN2(n634), .IN3(n1711), .Q(n1710));
   XOR2X1 U1468 (.IN1(n649), .IN2(n684), .Q(n1711));
   XOR3X1 U1470 (.IN1(n655), .IN2(n2213), .IN3(n1196), .Q(n1713));
   XOR2X1 U1471 (.IN1(n2207), .IN2(n2200), .Q(n1196));
   XOR2X1 U1472 (.IN1(n2221), .IN2(n638), .Q(n1195));
   XOR2X1 U1473 (.IN1(n1714), .IN2(n653), .Q(n1194));
   AOI22X1 U1474 (.IN1(n706), .IN2(block[30]), .IN3(new_block[30]), .IN4(n834), .QN(n1707)
          );
   OA22X1 U1475 (.IN1(new_block[30]), .IN2(n443), .IN3(block[30]), .IN4(n768), .Q(n1706)
          );
   AO221X1 U1476 (.IN1(n459), .IN2(new_sboxw[29]), .IN3(n144), .IN4(new_block[29]), .IN5(
          n1715), .Q(n2103));
   OAI222X1 U1477 (.IN1(n1716), .IN2(n2182), .IN3(round_key[29]), .IN4(n1717), .IN5(n1718)
          , .IN6(n971), .QN(n1715));
   XOR3X1 U1479 (.IN1(n667), .IN2(n651), .IN3(n1643), .Q(n1720));
   XOR2X1 U1480 (.IN1(n2183), .IN2(n649), .Q(n1643));
   XOR2X1 U1481 (.IN1(n2184), .IN2(new_block[28]), .Q(n1714));
   XOR3X1 U1483 (.IN1(n1207), .IN2(n2217), .IN3(n1208), .Q(n1721));
   XOR2X1 U1484 (.IN1(n666), .IN2(n2200), .Q(n1208));
   XNOR2X1 U1485 (.IN1(n695), .IN2(n742), .Q(n1223));
   XOR2X1 U1486 (.IN1(n2215), .IN2(n1237), .Q(n1207));
   XOR2X1 U1487 (.IN1(n707), .IN2(n638), .Q(n1237));
   XNOR2X1 U1488 (.IN1(n634), .IN2(n698), .Q(n1210));
   XOR2X1 U1489 (.IN1(n669), .IN2(n653), .Q(n1206));
   AOI22X1 U1490 (.IN1(n785), .IN2(block[29]), .IN3(new_block[29]), .IN4(n816), .QN(n1717)
          );
   OA22X1 U1491 (.IN1(new_block[29]), .IN2(n442), .IN3(block[29]), .IN4(n768), .Q(n1716)
          );
   AO221X1 U1492 (.IN1(n459), .IN2(new_sboxw[28]), .IN3(n144), .IN4(new_block[28]), .IN5(
          n1722), .Q(n2104));
   OAI222X1 U1493 (.IN1(n1723), .IN2(n2184), .IN3(round_key[28]), .IN4(n1724), .IN5(n1725)
          , .IN6(n971), .QN(n1722));
   XOR3X1 U1495 (.IN1(n633), .IN2(n667), .IN3(n1728), .Q(n1727));
   XOR2X1 U1496 (.IN1(n653), .IN2(n684), .Q(n1728));
   XOR2X1 U1497 (.IN1(n1241), .IN2(n740), .Q(n684));
   XOR2X1 U1498 (.IN1(n696), .IN2(n639), .Q(n653));
   XOR2X1 U1499 (.IN1(round_key[27]), .IN2(new_block[27]), .Q(n696));
   XNOR2X1 U1500 (.IN1(n169), .IN2(round_key[20]), .Q(n667));
   XNOR2X1 U1501 (.IN1(n184), .IN2(round_key[12]), .Q(n633));
   XOR3X1 U1503 (.IN1(n1220), .IN2(n2219), .IN3(n1221), .Q(n1729));
   XOR2X1 U1504 (.IN1(n666), .IN2(n1654), .Q(n1221));
   XOR2X1 U1505 (.IN1(n651), .IN2(n1730), .Q(n1654));
   XOR2X1 U1506 (.IN1(n2203), .IN2(n2199), .Q(n666));
   XNOR2X1 U1507 (.IN1(n710), .IN2(n742), .Q(n1239));
   XNOR2X1 U1508 (.IN1(n197), .IN2(round_key[4]), .Q(n1184));
   XOR2X1 U1509 (.IN1(n2217), .IN2(n1663), .Q(n1220));
   XNOR2X1 U1510 (.IN1(n723), .IN2(n2215), .Q(n1663));
   XNOR2X1 U1511 (.IN1(n649), .IN2(n1662), .Q(n1224));
   XOR2X1 U1512 (.IN1(n714), .IN2(n634), .Q(n1662));
   XOR2X1 U1513 (.IN1(n669), .IN2(n1653), .Q(n1219));
   XOR2X1 U1514 (.IN1(n2181), .IN2(n1731), .Q(n1653));
   XNOR2X1 U1515 (.IN1(n656), .IN2(n1665), .Q(n669));
   AOI22X1 U1516 (.IN1(n679), .IN2(block[28]), .IN3(new_block[28]), .IN4(n800), .QN(n1724)
          );
   OA22X1 U1517 (.IN1(new_block[28]), .IN2(n446), .IN3(block[28]), .IN4(n768), .Q(n1723)
          );
   AO221X1 U1518 (.IN1(n459), .IN2(new_sboxw[27]), .IN3(n144), .IN4(new_block[27]), .IN5(
          n1732), .Q(n2105));
   OAI222X1 U1519 (.IN1(n1733), .IN2(n2185), .IN3(round_key[27]), .IN4(n1734), .IN5(n1735)
          , .IN6(n939), .QN(n1732));
   XOR2X1 U1520 (.IN1(n1736), .IN2(n1737), .Q(n1735));
   XOR2X1 U1523 (.IN1(n1253), .IN2(n740), .Q(n698));
   XOR2X1 U1524 (.IN1(n711), .IN2(n639), .Q(n1665));
   XOR2X1 U1525 (.IN1(round_key[26]), .IN2(new_block[26]), .Q(n711));
   XOR2X1 U1526 (.IN1(n170), .IN2(n2193), .Q(n1241));
   XOR2X1 U1527 (.IN1(n185), .IN2(n2208), .Q(n695));
   XOR3X1 U1528 (.IN1(n1233), .IN2(n1240), .IN3(n1739), .Q(n1736));
   XOR3X1 U1529 (.IN1(n1234), .IN2(n2221), .IN3(n1235), .Q(n1739));
   XNOR2X1 U1530 (.IN1(n1667), .IN2(n1730), .Q(n1235));
   XNOR2X1 U1531 (.IN1(n713), .IN2(n2203), .Q(n1730));
   XOR2X1 U1532 (.IN1(n2205), .IN2(n1268), .Q(n1667));
   XNOR2X1 U1533 (.IN1(n199), .IN2(round_key[3]), .Q(n1236));
   XOR2X1 U1534 (.IN1(n2217), .IN2(n1266), .Q(n1234));
   XOR2X1 U1535 (.IN1(n737), .IN2(n638), .Q(n1266));
   XNOR2X1 U1536 (.IN1(n649), .IN2(n728), .Q(n1240));
   XOR2X1 U1538 (.IN1(n726), .IN2(n656), .Q(n1731));
   XOR2X1 U1539 (.IN1(n1712), .IN2(n1685), .Q(n1666));
   AOI22X1 U1540 (.IN1(n664), .IN2(block[27]), .IN3(new_block[27]), .IN4(n833), .QN(n1734)
          );
   OA22X1 U1541 (.IN1(new_block[27]), .IN2(n897), .IN3(block[27]), .IN4(n768), .Q(n1733)
          );
   AO221X1 U1542 (.IN1(n459), .IN2(new_sboxw[26]), .IN3(n144), .IN4(new_block[26]), .IN5(
          n1740), .Q(n2106));
   OAI222X1 U1543 (.IN1(n1741), .IN2(n2186), .IN3(round_key[26]), .IN4(n1742), .IN5(n1743)
          , .IN6(n939), .QN(n1740));
   XOR3X1 U1545 (.IN1(n710), .IN2(n1253), .IN3(n1746), .Q(n1745));
   XOR2X1 U1546 (.IN1(n726), .IN2(n714), .Q(n1746));
   XOR2X1 U1547 (.IN1(round_key[25]), .IN2(new_block[25]), .Q(n726));
   XOR2X1 U1548 (.IN1(n171), .IN2(n2194), .Q(n1253));
   XOR2X1 U1549 (.IN1(n186), .IN2(n2209), .Q(n710));
   XOR3X1 U1551 (.IN1(n707), .IN2(n1250), .IN3(n1252), .Q(n1747));
   XOR2X1 U1552 (.IN1(n1268), .IN2(n635), .Q(n1252));
   XNOR2X1 U1553 (.IN1(n744), .IN2(n742), .Q(n1268));
   XOR2X1 U1554 (.IN1(n655), .IN2(n638), .Q(n1250));
   XOR2X1 U1555 (.IN1(new_block[7]), .IN2(round_key[7]), .Q(n638));
   XOR2X1 U1556 (.IN1(n200), .IN2(n2222), .Q(n707));
   XNOR2X1 U1557 (.IN1(n1685), .IN2(n1676), .Q(n1251));
   XOR2X1 U1558 (.IN1(n740), .IN2(n634), .Q(n1255));
   AOI22X1 U1559 (.IN1(n697), .IN2(block[26]), .IN3(new_block[26]), .IN4(n437), .QN(n1742)
          );
   OA22X1 U1560 (.IN1(new_block[26]), .IN2(n850), .IN3(block[26]), .IN4(n768), .Q(n1741)
          );
   AO221X1 U1561 (.IN1(n459), .IN2(new_sboxw[25]), .IN3(n144), .IN4(new_block[25]), .IN5(
          n1748), .Q(n2107));
   OAI222X1 U1562 (.IN1(n1749), .IN2(n2187), .IN3(round_key[25]), .IN4(n1750), .IN5(n1751)
          , .IN6(n939), .QN(n1748));
   XOR3X1 U1564 (.IN1(n713), .IN2(n714), .IN3(n1754), .Q(n1753));
   XNOR2X1 U1565 (.IN1(n1685), .IN2(n728), .Q(n1754));
   XOR2X1 U1566 (.IN1(n1279), .IN2(n740), .Q(n728));
   XNOR2X1 U1567 (.IN1(n743), .IN2(n639), .Q(n1685));
   XOR2X1 U1568 (.IN1(round_key[24]), .IN2(new_block[24]), .Q(n743));
   XOR2X1 U1569 (.IN1(n172), .IN2(n2195), .Q(n714));
   XOR2X1 U1570 (.IN1(n187), .IN2(n2210), .Q(n713));
   XOR3X1 U1572 (.IN1(n723), .IN2(n738), .IN3(n1265), .Q(n1755));
   XOR2X1 U1573 (.IN1(n2202), .IN2(n635), .Q(n1265));
   XOR2X1 U1574 (.IN1(n648), .IN2(n742), .Q(n635));
   XOR2X1 U1575 (.IN1(new_block[15]), .IN2(round_key[15]), .Q(n742));
   XOR2X1 U1576 (.IN1(n2215), .IN2(n2217), .Q(n738));
   XNOR2X1 U1577 (.IN1(n193), .IN2(round_key[6]), .Q(n655));
   XOR2X1 U1578 (.IN1(n201), .IN2(n2223), .Q(n723));
   XNOR2X1 U1579 (.IN1(n1277), .IN2(n1676), .Q(n1264));
   XOR2X1 U1580 (.IN1(n656), .IN2(n639), .Q(n1676));
   XOR2X1 U1581 (.IN1(n634), .IN2(n649), .Q(n739));
   AOI22X1 U1583 (.IN1(n664), .IN2(block[25]), .IN3(new_block[25]), .IN4(n833), .QN(n1750)
          );
   OA22X1 U1584 (.IN1(new_block[25]), .IN2(n868), .IN3(block[25]), .IN4(n768), .Q(n1749)
          );
   AO221X1 U1585 (.IN1(n459), .IN2(new_sboxw[24]), .IN3(n144), .IN4(new_block[24]), .IN5(
          n1756), .Q(n2108));
   OAI222X1 U1586 (.IN1(n1757), .IN2(n2188), .IN3(round_key[24]), .IN4(n1758), .IN5(n1759)
          , .IN6(n939), .QN(n1756));
   XOR3X1 U1588 (.IN1(n740), .IN2(n744), .IN3(n1762), .Q(n1761));
   XOR2X1 U1589 (.IN1(n649), .IN2(n639), .Q(n1762));
   XOR2X1 U1590 (.IN1(round_key[31]), .IN2(new_block[31]), .Q(n639));
   XOR2X1 U1592 (.IN1(n188), .IN2(n2211), .Q(n744));
   XOR3X1 U1595 (.IN1(n671), .IN2(n737), .IN3(n2202), .Q(n1763));
   XNOR2X1 U1596 (.IN1(n2203), .IN2(n651), .Q(n1278));
   XNOR2X1 U1597 (.IN1(n182), .IN2(round_key[13]), .Q(n651));
   XNOR2X1 U1598 (.IN1(n180), .IN2(round_key[14]), .Q(n648));
   XOR2X1 U1599 (.IN1(n202), .IN2(n2224), .Q(n737));
   XNOR2X1 U1600 (.IN1(n195), .IN2(round_key[5]), .Q(n671));
   XOR2X1 U1601 (.IN1(n656), .IN2(n1712), .Q(n1277));
   XOR2X1 U1602 (.IN1(n2182), .IN2(new_block[29]), .Q(n1712));
   XNOR2X1 U1603 (.IN1(n2180), .IN2(new_block[30]), .Q(n656));
   XOR2X1 U1604 (.IN1(n173), .IN2(n2196), .Q(n1279));
   AOI22X1 U1605 (.IN1(n697), .IN2(block[24]), .IN3(new_block[24]), .IN4(n816), .QN(n1758)
          );
   OA22X1 U1606 (.IN1(new_block[24]), .IN2(n443), .IN3(block[24]), .IN4(n753), .Q(n1757)
          );
   AO221X1 U1607 (.IN1(n459), .IN2(new_sboxw[23]), .IN3(n664), .IN4(n1765), .IN5(n1766), .
          Q(n2109));
   OAI222X1 U1608 (.IN1(n1767), .IN2(n164), .IN3(n2189), .IN4(n1768), .IN5(n1769), .IN6(
          n939), .QN(n1766));
   XOR2X1 U1611 (.IN1(n2149), .IN2(n791), .Q(n1290));
   XOR2X1 U1612 (.IN1(n755), .IN2(n767), .Q(n1289));
   XOR2X1 U1614 (.IN1(n758), .IN2(n790), .Q(n1773));
   XOR2X1 U1616 (.IN1(round_key[55]), .IN2(block[55]), .Q(n1765));
   AO221X1 U1617 (.IN1(n459), .IN2(new_sboxw[22]), .IN3(n785), .IN4(n1774), .IN5(n1775), .
          Q(n2110));
   OAI222X1 U1618 (.IN1(n1776), .IN2(n166), .IN3(n2190), .IN4(n1777), .IN5(n1778), .IN6(
          n939), .QN(n1775));
   XOR3X1 U1620 (.IN1(n1300), .IN2(n2169), .IN3(n1301), .Q(n1781));
   XOR2X1 U1621 (.IN1(n2149), .IN2(n776), .Q(n1301));
   XOR2X1 U1622 (.IN1(n2173), .IN2(n2167), .Q(n1300));
   XOR3X1 U1623 (.IN1(n758), .IN2(n771), .IN3(n1782), .Q(n1780));
   XOR2X1 U1624 (.IN1(n806), .IN2(n1303), .Q(n1782));
   XOR2X1 U1625 (.IN1(n825), .IN2(n760), .Q(n1303));
   XOR2X1 U1627 (.IN1(round_key[54]), .IN2(block[54]), .Q(n1774));
   AO221X1 U1628 (.IN1(n459), .IN2(new_sboxw[21]), .IN3(n736), .IN4(n1783), .IN5(n1784), .
          Q(n2111));
   OAI222X1 U1629 (.IN1(n1785), .IN2(n167), .IN3(n2191), .IN4(n1786), .IN5(n1787), .IN6(
          n939), .QN(n1784));
   XOR3X1 U1631 (.IN1(n1312), .IN2(n2171), .IN3(n1313), .Q(n1790));
   XNOR2X1 U1632 (.IN1(n792), .IN2(n776), .Q(n1313));
   XOR2X1 U1633 (.IN1(n788), .IN2(n2167), .Q(n1312));
   XOR2X1 U1634 (.IN1(n2175), .IN2(n750), .Q(n772));
   XOR3X1 U1635 (.IN1(n1926), .IN2(n809), .IN3(n759), .Q(n1789));
   XOR2X1 U1636 (.IN1(n771), .IN2(n790), .Q(n759));
   XNOR2X1 U1637 (.IN1(n215), .IN2(round_key[52]), .Q(n809));
   XNOR2X1 U1639 (.IN1(n777), .IN2(n1340), .Q(n1316));
   XOR2X1 U1640 (.IN1(n840), .IN2(n760), .Q(n1340));
   XOR2X1 U1641 (.IN1(n2159), .IN2(n2156), .Q(n1315));
   XOR2X1 U1642 (.IN1(round_key[53]), .IN2(block[53]), .Q(n1783));
   AO221X1 U1643 (.IN1(n459), .IN2(new_sboxw[20]), .IN3(n727), .IN4(n1792), .IN5(n1793), .
          Q(n2112));
   OAI222X1 U1644 (.IN1(n1794), .IN2(n169), .IN3(n2192), .IN4(n1795), .IN5(n1796), .IN6(
          n939), .QN(n1793));
   XOR3X1 U1645 (.IN1(n1322), .IN2(n1797), .IN3(n1798), .Q(n1796));
   XOR3X1 U1646 (.IN1(n1325), .IN2(n2173), .IN3(n1326), .Q(n1798));
   XNOR2X1 U1647 (.IN1(n792), .IN2(n803), .Q(n1326));
   XNOR2X1 U1648 (.IN1(n2147), .IN2(n1799), .Q(n803));
   XNOR2X1 U1649 (.IN1(n2145), .IN2(n1419), .Q(n792));
   XNOR2X1 U1650 (.IN1(n241), .IN2(round_key[36]), .Q(n755));
   XNOR2X1 U1651 (.IN1(n788), .IN2(n807), .Q(n1325));
   XNOR2X1 U1652 (.IN1(n767), .IN2(n1800), .Q(n807));
   XOR2X1 U1653 (.IN1(n2169), .IN2(n822), .Q(n788));
   XOR2X1 U1654 (.IN1(n838), .IN2(n750), .Q(n822));
   XNOR2X1 U1657 (.IN1(n826), .IN2(n2143), .Q(n776));
   XOR2X1 U1658 (.IN1(n216), .IN2(n2150), .Q(n826));
   XOR2X1 U1659 (.IN1(n1338), .IN2(n875), .Q(n806));
   XNOR2X1 U1660 (.IN1(n1943), .IN2(new_block[60]), .Q(n808));
   XNOR2X1 U1661 (.IN1(n229), .IN2(round_key[44]), .Q(n790));
   XOR2X1 U1662 (.IN1(n1411), .IN2(n1410), .Q(n1322));
   XOR2X1 U1663 (.IN1(n771), .IN2(n1424), .Q(n1410));
   XNOR2X1 U1664 (.IN1(n843), .IN2(n2159), .Q(n1424));
   XOR2X1 U1665 (.IN1(n1926), .IN2(n1422), .Q(n1411));
   XNOR2X1 U1666 (.IN1(n857), .IN2(n777), .Q(n1422));
   XOR2X1 U1667 (.IN1(round_key[52]), .IN2(block[52]), .Q(n1792));
   AO221X1 U1668 (.IN1(n460), .IN2(new_sboxw[19]), .IN3(n736), .IN4(n1802), .IN5(n1803), .
          Q(n2113));
   OAI222X1 U1669 (.IN1(n1804), .IN2(n170), .IN3(n2193), .IN4(n1805), .IN5(n1806), .IN6(
          n939), .QN(n1803));
   XOR3X1 U1670 (.IN1(n1333), .IN2(n1807), .IN3(n1808), .Q(n1806));
   XOR3X1 U1671 (.IN1(n1336), .IN2(n2175), .IN3(n1337), .Q(n1808));
   XOR2X1 U1672 (.IN1(n820), .IN2(n1799), .Q(n1337));
   XNOR2X1 U1673 (.IN1(n858), .IN2(n2145), .Q(n1799));
   XOR2X1 U1674 (.IN1(n2147), .IN2(n1442), .Q(n820));
   XNOR2X1 U1675 (.IN1(n243), .IN2(round_key[35]), .Q(n821));
   XOR2X1 U1676 (.IN1(n824), .IN2(n1800), .Q(n1336));
   XNOR2X1 U1677 (.IN1(n839), .IN2(n2169), .Q(n1800));
   XOR2X1 U1678 (.IN1(n767), .IN2(n856), .Q(n824));
   XNOR2X1 U1681 (.IN1(n841), .IN2(n2143), .Q(n1419));
   XOR2X1 U1682 (.IN1(n217), .IN2(n2151), .Q(n841));
   XOR2X1 U1683 (.IN1(n1351), .IN2(n875), .Q(n1791));
   XOR2X1 U1684 (.IN1(round_key[59]), .IN2(new_block[59]), .Q(n825));
   XOR2X1 U1685 (.IN1(n230), .IN2(n2162), .Q(n1338));
   XOR2X1 U1686 (.IN1(n1421), .IN2(n1423), .Q(n1333));
   XOR2X1 U1688 (.IN1(n1810), .IN2(n1364), .Q(n1421));
   XNOR2X1 U1689 (.IN1(n873), .IN2(n760), .Q(n1364));
   XOR2X1 U1690 (.IN1(round_key[51]), .IN2(block[51]), .Q(n1802));
   AO221X1 U1691 (.IN1(n460), .IN2(new_sboxw[18]), .IN3(n631), .IN4(n1811), .IN5(n1812), .
          Q(n2114));
   OAI222X1 U1692 (.IN1(n1813), .IN2(n171), .IN3(n2194), .IN4(n1814), .IN5(n1815), .IN6(
          n939), .QN(n1812));
   XNOR2X1 U1695 (.IN1(n1442), .IN2(n836), .Q(n1350));
   XNOR2X1 U1696 (.IN1(n856), .IN2(n844), .Q(n1349));
   XNOR2X1 U1697 (.IN1(n872), .IN2(n750), .Q(n856));
   XOR2X1 U1698 (.IN1(n244), .IN2(n2176), .Q(n838));
   XOR3X1 U1699 (.IN1(n1351), .IN2(n840), .IN3(n1818), .Q(n1816));
   XOR2X1 U1700 (.IN1(n843), .IN2(n858), .Q(n1818));
   XOR2X1 U1701 (.IN1(n218), .IN2(n2152), .Q(n858));
   XOR2X1 U1702 (.IN1(round_key[58]), .IN2(new_block[58]), .Q(n840));
   XOR2X1 U1703 (.IN1(n231), .IN2(n2163), .Q(n1351));
   XOR2X1 U1704 (.IN1(n1434), .IN2(n1433), .Q(n1346));
   XOR2X1 U1705 (.IN1(n875), .IN2(n758), .Q(n1433));
   XOR2X1 U1706 (.IN1(n1912), .IN2(n760), .Q(n1434));
   XOR2X1 U1707 (.IN1(round_key[63]), .IN2(new_block[63]), .Q(n760));
   XOR2X1 U1708 (.IN1(round_key[50]), .IN2(block[50]), .Q(n1811));
   AO221X1 U1709 (.IN1(n460), .IN2(new_sboxw[17]), .IN3(n706), .IN4(n1819), .IN5(n1820), .
          Q(n2115));
   OAI222X1 U1710 (.IN1(n1821), .IN2(n172), .IN3(n2195), .IN4(n1822), .IN5(n1823), .IN6(
          n939), .QN(n1820));
   XOR3X1 U1711 (.IN1(n1358), .IN2(n1824), .IN3(n1825), .Q(n1823));
   XOR3X1 U1712 (.IN1(n839), .IN2(n1361), .IN3(n1362), .Q(n1825));
   XNOR2X1 U1713 (.IN1(n854), .IN2(n836), .Q(n1362));
   XOR2X1 U1714 (.IN1(n2145), .IN2(n2143), .Q(n836));
   XOR2X1 U1715 (.IN1(n861), .IN2(n844), .Q(n1361));
   XOR2X1 U1716 (.IN1(n751), .IN2(n750), .Q(n844));
   XOR2X1 U1717 (.IN1(new_block[39]), .IN2(round_key[39]), .Q(n750));
   XOR2X1 U1718 (.IN1(n245), .IN2(n2177), .Q(n839));
   XOR2X1 U1721 (.IN1(n870), .IN2(n756), .Q(n1442));
   XOR2X1 U1722 (.IN1(n219), .IN2(n2153), .Q(n870));
   XOR2X1 U1723 (.IN1(n1373), .IN2(n875), .Q(n860));
   XOR2X1 U1724 (.IN1(n232), .IN2(n2164), .Q(n843));
   XOR2X1 U1725 (.IN1(round_key[57]), .IN2(new_block[57]), .Q(n857));
   XOR2X1 U1726 (.IN1(n871), .IN2(n1452), .Q(n1358));
   XNOR2X1 U1727 (.IN1(n2159), .IN2(n771), .Q(n1452));
   XNOR2X1 U1728 (.IN1(n225), .IN2(round_key[46]), .Q(n758));
   XOR2X1 U1729 (.IN1(n777), .IN2(n1810), .Q(n871));
   XOR2X1 U1730 (.IN1(n1919), .IN2(new_block[62]), .Q(n777));
   XOR2X1 U1731 (.IN1(round_key[49]), .IN2(block[49]), .Q(n1819));
   AO221X1 U1732 (.IN1(n460), .IN2(new_sboxw[16]), .IN3(n727), .IN4(n1827), .IN5(n1828), .
          Q(n2116));
   OAI222X1 U1733 (.IN1(n1829), .IN2(n173), .IN3(n2196), .IN4(n1830), .IN5(n1831), .IN6(
          n939), .QN(n1828));
   XOR2X1 U1736 (.IN1(n2145), .IN2(n2147), .Q(n854));
   XNOR2X1 U1737 (.IN1(n213), .IN2(round_key[53]), .Q(n791));
   XNOR2X1 U1738 (.IN1(n211), .IN2(round_key[54]), .Q(n775));
   XOR2X1 U1739 (.IN1(n2169), .IN2(n2171), .Q(n861));
   XNOR2X1 U1740 (.IN1(n239), .IN2(round_key[37]), .Q(n767));
   XNOR2X1 U1741 (.IN1(n237), .IN2(round_key[38]), .Q(n751));
   XOR2X1 U1742 (.IN1(n246), .IN2(n2178), .Q(n872));
   XOR3X1 U1743 (.IN1(n1926), .IN2(n875), .IN3(n1835), .Q(n1833));
   XOR2X1 U1744 (.IN1(n756), .IN2(n771), .Q(n1835));
   XNOR2X1 U1745 (.IN1(n227), .IN2(round_key[45]), .Q(n771));
   XNOR2X1 U1746 (.IN1(n209), .IN2(round_key[55]), .Q(n756));
   XNOR2X1 U1747 (.IN1(n222), .IN2(round_key[47]), .Q(n875));
   XOR2X1 U1748 (.IN1(n1935), .IN2(new_block[61]), .Q(n1810));
   XOR2X1 U1749 (.IN1(n873), .IN2(n1373), .Q(n1832));
   XOR2X1 U1750 (.IN1(n233), .IN2(n2165), .Q(n1373));
   XOR2X1 U1751 (.IN1(round_key[56]), .IN2(new_block[56]), .Q(n873));
   XOR2X1 U1752 (.IN1(round_key[48]), .IN2(block[48]), .Q(n1827));
   AO221X1 U1753 (.IN1(n460), .IN2(new_sboxw[15]), .IN3(n631), .IN4(n1836), .IN5(n1837), .
          Q(n2117));
   OAI222X1 U1754 (.IN1(n1838), .IN2(n177), .IN3(n2197), .IN4(n1839), .IN5(n1840), .IN6(
          n939), .QN(n1837));
   XOR3X1 U1756 (.IN1(n990), .IN2(n987), .IN3(n991), .Q(n1843));
   XOR2X1 U1757 (.IN1(n1809), .IN2(n1011), .Q(n991));
   XOR2X1 U1758 (.IN1(n1634), .IN2(n1623), .Q(n987));
   XOR3X1 U1760 (.IN1(n888), .IN2(n899), .IN3(n1844), .Q(n1841));
   XOR2X1 U1761 (.IN1(n886), .IN2(n930), .Q(n1844));
   XOR2X1 U1762 (.IN1(round_key[79]), .IN2(block[79]), .Q(n1836));
   AO221X1 U1763 (.IN1(n460), .IN2(new_sboxw[14]), .IN3(n646), .IN4(n1845), .IN5(n1846), .
          Q(n2118));
   OAI222X1 U1764 (.IN1(n1847), .IN2(n180), .IN3(n2201), .IN4(n1848), .IN5(n1849), .IN6(
          n939), .QN(n1846));
   XOR2X1 U1767 (.IN1(n1809), .IN2(n1764), .Q(n1003));
   XOR2X1 U1768 (.IN1(n1854), .IN2(n1613), .Q(n1000));
   XOR2X1 U1769 (.IN1(n890), .IN2(n905), .Q(n1851));
   XOR3X1 U1770 (.IN1(n1614), .IN2(n901), .IN3(n1855), .Q(n1850));
   XOR2X1 U1771 (.IN1(n999), .IN2(n929), .Q(n1855));
   XOR2X1 U1772 (.IN1(n946), .IN2(n886), .Q(n999));
   XOR2X1 U1773 (.IN1(round_key[78]), .IN2(block[78]), .Q(n1845));
   AO221X1 U1774 (.IN1(n460), .IN2(new_sboxw[13]), .IN3(n631), .IN4(n1856), .IN5(n1857), .
          Q(n2119));
   OAI222X1 U1775 (.IN1(n1858), .IN2(n182), .IN3(n2204), .IN4(n1859), .IN5(n1860), .IN6(
          n939), .QN(n1857));
   XOR2X1 U1778 (.IN1(n1479), .IN2(n1853), .Q(n1016));
   XOR2X1 U1779 (.IN1(n1870), .IN2(n941), .Q(n1015));
   XOR2X1 U1780 (.IN1(n1480), .IN2(n1613), .Q(n1012));
   XNOR2X1 U1781 (.IN1(n944), .IN2(n888), .Q(n903));
   XOR2X1 U1784 (.IN1(n1693), .IN2(n1036), .Q(n1013));
   XOR2X1 U1785 (.IN1(n962), .IN2(n886), .Q(n1036));
   XOR2X1 U1786 (.IN1(n884), .IN2(n917), .Q(n1864));
   XNOR2X1 U1787 (.IN1(n274), .IN2(round_key[76]), .Q(n884));
   XOR2X1 U1788 (.IN1(round_key[77]), .IN2(block[77]), .Q(n1856));
   AO221X1 U1789 (.IN1(n460), .IN2(new_sboxw[12]), .IN3(n646), .IN4(n1865), .IN5(n1866), .
          Q(n2120));
   OAI222X1 U1790 (.IN1(n1867), .IN2(n184), .IN3(n2206), .IN4(n1868), .IN5(n1869), .IN6(
          n926), .QN(n1866));
   XNOR2X1 U1793 (.IN1(n1479), .IN2(n1490), .Q(n1028));
   XOR2X1 U1794 (.IN1(n1011), .IN2(n1873), .Q(n1490));
   XOR2X1 U1795 (.IN1(n1772), .IN2(n1501), .Q(n1479));
   XOR2X1 U1796 (.IN1(n1872), .IN2(n1499), .Q(n1027));
   XNOR2X1 U1797 (.IN1(n956), .IN2(n1870), .Q(n1499));
   XOR2X1 U1798 (.IN1(n1480), .IN2(n1489), .Q(n1024));
   XOR2X1 U1799 (.IN1(n1623), .IN2(n1874), .Q(n1489));
   XOR2X1 U1800 (.IN1(n1875), .IN2(n947), .Q(n1480));
   XOR2X1 U1801 (.IN1(n959), .IN2(n888), .Q(n947));
   XOR2X1 U1803 (.IN1(n1041), .IN2(n990), .Q(n929));
   XNOR2X1 U1804 (.IN1(n288), .IN2(round_key[68]), .Q(n989));
   XOR2X1 U1806 (.IN1(n1703), .IN2(n1498), .Q(n1025));
   XNOR2X1 U1807 (.IN1(n977), .IN2(n1693), .Q(n1498));
   XNOR2X1 U1808 (.IN1(n943), .IN2(n883), .Q(n1853));
   XOR2X1 U1809 (.IN1(n275), .IN2(n1817), .Q(n943));
   XOR2X1 U1810 (.IN1(n930), .IN2(n1634), .Q(n1876));
   XOR2X1 U1811 (.IN1(n1642), .IN2(new_block[92]), .Q(n1854));
   XNOR2X1 U1812 (.IN1(n260), .IN2(round_key[84]), .Q(n930));
   XOR2X1 U1813 (.IN1(round_key[76]), .IN2(block[76]), .Q(n1865));
   AO221X1 U1814 (.IN1(n460), .IN2(new_sboxw[11]), .IN3(n679), .IN4(n1877), .IN5(n1878), .
          Q(n2121));
   OAI222X1 U1815 (.IN1(n1879), .IN2(n185), .IN3(n2208), .IN4(n1880), .IN5(n1881), .IN6(
          n926), .QN(n1878));
   XOR3X1 U1817 (.IN1(n1037), .IN2(n1040), .IN3(n1042), .Q(n1884));
   XNOR2X1 U1818 (.IN1(n1503), .IN2(n1873), .Q(n1042));
   XNOR2X1 U1819 (.IN1(n975), .IN2(n1772), .Q(n1873));
   XOR2X1 U1820 (.IN1(n1788), .IN2(n1522), .Q(n1503));
   XOR2X1 U1821 (.IN1(n1872), .IN2(n972), .Q(n1040));
   XNOR2X1 U1823 (.IN1(n963), .IN2(n1875), .Q(n1874));
   XOR2X1 U1824 (.IN1(n1001), .IN2(n978), .Q(n1502));
   XOR2X1 U1826 (.IN1(n1053), .IN2(n990), .Q(n941));
   XOR2X1 U1827 (.IN1(n289), .IN2(n1900), .Q(n1041));
   XOR3X1 U1828 (.IN1(n1885), .IN2(n1501), .IN3(n1038), .Q(n1882));
   XOR2X1 U1829 (.IN1(n1703), .IN2(n1063), .Q(n1038));
   XOR2X1 U1830 (.IN1(n1077), .IN2(n886), .Q(n1063));
   XNOR2X1 U1831 (.IN1(n960), .IN2(n883), .Q(n1501));
   XOR2X1 U1832 (.IN1(n276), .IN2(n1826), .Q(n960));
   XOR2X1 U1833 (.IN1(n944), .IN2(n946), .Q(n1885));
   XOR2X1 U1834 (.IN1(n261), .IN2(n1719), .Q(n946));
   XOR2X1 U1835 (.IN1(round_key[91]), .IN2(new_block[91]), .Q(n944));
   XOR2X1 U1836 (.IN1(round_key[75]), .IN2(block[75]), .Q(n1877));
   AO221X1 U1837 (.IN1(n460), .IN2(new_sboxw[10]), .IN3(n736), .IN4(n1886), .IN5(n1887), .
          Q(n2122));
   OAI222X1 U1838 (.IN1(n1888), .IN2(n186), .IN3(n2209), .IN4(n1889), .IN5(n1890), .IN6(
          n926), .QN(n1887));
   XOR3X1 U1840 (.IN1(n1054), .IN2(n1051), .IN3(n1055), .Q(n1893));
   XOR2X1 U1841 (.IN1(n1522), .IN2(n1513), .Q(n1055));
   XNOR2X1 U1842 (.IN1(n978), .IN2(n1512), .Q(n1051));
   XNOR2X1 U1843 (.IN1(n1531), .IN2(n888), .Q(n978));
   XOR2X1 U1844 (.IN1(n990), .IN2(n890), .Q(n1054));
   XOR2X1 U1846 (.IN1(n290), .IN2(n1901), .Q(n1053));
   XOR3X1 U1847 (.IN1(n959), .IN2(n962), .IN3(n1894), .Q(n1891));
   XOR2X1 U1848 (.IN1(n975), .IN2(n1050), .Q(n1894));
   XOR2X1 U1849 (.IN1(n901), .IN2(n886), .Q(n1050));
   XOR2X1 U1850 (.IN1(new_block[87]), .IN2(round_key[87]), .Q(n886));
   XOR2X1 U1851 (.IN1(n277), .IN2(n1834), .Q(n975));
   XOR2X1 U1852 (.IN1(n262), .IN2(n1726), .Q(n962));
   XOR2X1 U1853 (.IN1(round_key[90]), .IN2(new_block[90]), .Q(n959));
   XOR2X1 U1854 (.IN1(round_key[74]), .IN2(block[74]), .Q(n1886));
   AO221X1 U1855 (.IN1(n460), .IN2(new_sboxw[9]), .IN3(n706), .IN4(n1895), .IN5(n1896), .Q(
          n2123));
   OAI222X1 U1856 (.IN1(n1897), .IN2(n187), .IN3(n2210), .IN4(n1898), .IN5(n1899), .IN6(
          n926), .QN(n1896));
   XOR2X1 U1859 (.IN1(n1771), .IN2(n1513), .Q(n1068));
   XOR2X1 U1860 (.IN1(n899), .IN2(n883), .Q(n1513));
   XNOR2X1 U1861 (.IN1(n1078), .IN2(n1512), .Q(n1065));
   XOR2X1 U1862 (.IN1(n1614), .IN2(n888), .Q(n1512));
   XOR2X1 U1864 (.IN1(n1080), .IN2(n990), .Q(n972));
   XOR2X1 U1865 (.IN1(n291), .IN2(n1902), .Q(n956));
   XNOR2X1 U1867 (.IN1(n1522), .IN2(n1064), .Q(n1904));
   XNOR2X1 U1868 (.IN1(n1075), .IN2(n883), .Q(n1522));
   XOR2X1 U1869 (.IN1(n263), .IN2(n1738), .Q(n977));
   XOR2X1 U1870 (.IN1(round_key[89]), .IN2(new_block[89]), .Q(n963));
   XOR2X1 U1871 (.IN1(round_key[73]), .IN2(block[73]), .Q(n1895));
   AO221X1 U1872 (.IN1(n460), .IN2(new_sboxw[8]), .IN3(n727), .IN4(n1905), .IN5(n1906), .Q(
          n2124));
   OAI222X1 U1873 (.IN1(n1907), .IN2(n188), .IN3(n2211), .IN4(n1908), .IN5(n1909), .IN6(
          n926), .QN(n1906));
   XNOR2X1 U1876 (.IN1(n1772), .IN2(n1011), .Q(n1903));
   XNOR2X1 U1877 (.IN1(n270), .IN2(round_key[78]), .Q(n899));
   XOR2X1 U1878 (.IN1(n1614), .IN2(n1001), .Q(n1078));
   XOR2X1 U1879 (.IN1(n1615), .IN2(new_block[94]), .Q(n1875));
   XOR2X1 U1880 (.IN1(n292), .IN2(n1910), .Q(n1080));
   XOR2X1 U1883 (.IN1(n883), .IN2(n917), .Q(n1913));
   XOR2X1 U1884 (.IN1(new_block[79]), .IN2(round_key[79]), .Q(n883));
   XOR2X1 U1885 (.IN1(round_key[72]), .IN2(block[72]), .Q(n1905));
   AO221X1 U1886 (.IN1(n461), .IN2(new_sboxw[7]), .IN3(n736), .IN4(n1914), .IN5(n1915), .Q(
          n2125));
   OAI222X1 U1887 (.IN1(n1916), .IN2(n190), .IN3(n2212), .IN4(n1917), .IN5(n1918), .IN6(
          n926), .QN(n1915));
   XOR3X1 U1889 (.IN1(n1541), .IN2(n1090), .IN3(n1091), .Q(n1920));
   XOR2X1 U1890 (.IN1(n1370), .IN2(n542), .Q(n1091));
   XOR2X1 U1891 (.IN1(n517), .IN2(n547), .Q(n1090));
   XOR2X1 U1893 (.IN1(n511), .IN2(n555), .Q(n1092));
   XOR2X1 U1894 (.IN1(round_key[103]), .IN2(block[103]), .Q(n1914));
   AO221X1 U1895 (.IN1(n461), .IN2(new_sboxw[6]), .IN3(n646), .IN4(n1921), .IN5(n1922), .Q(
          n2126));
   OAI222X1 U1896 (.IN1(n1923), .IN2(n193), .IN3(n2214), .IN4(n1924), .IN5(n1925), .IN6(
          n926), .QN(n1922));
   XOR3X1 U1898 (.IN1(n1102), .IN2(n1539), .IN3(n1103), .Q(n1928));
   XOR2X1 U1899 (.IN1(n1370), .IN2(n532), .Q(n1103));
   XOR2X1 U1900 (.IN1(n1549), .IN2(n531), .Q(n1102));
   XOR3X1 U1901 (.IN1(n1247), .IN2(n1093), .IN3(n527), .Q(n1927));
   XOR2X1 U1902 (.IN1(n509), .IN2(n1261), .Q(n527));
   XNOR2X1 U1904 (.IN1(n569), .IN2(n511), .Q(n1562));
   XOR2X1 U1905 (.IN1(round_key[102]), .IN2(block[102]), .Q(n1921));
   AO221X1 U1906 (.IN1(n461), .IN2(new_sboxw[5]), .IN3(n727), .IN4(n1929), .IN5(n1930), .Q(
          n2127));
   OAI222X1 U1907 (.IN1(n1931), .IN2(n195), .IN3(n2216), .IN4(n1932), .IN5(n1933), .IN6(
          n926), .QN(n1930));
   XOR2X1 U1910 (.IN1(n548), .IN2(n532), .Q(n1114));
   XOR2X1 U1911 (.IN1(n570), .IN2(n508), .Q(n532));
   XNOR2X1 U1912 (.IN1(n330), .IN2(round_key[100]), .Q(n517));
   XNOR2X1 U1913 (.IN1(n546), .IN2(n531), .Q(n1113));
   XOR3X1 U1914 (.IN1(n540), .IN2(n542), .IN3(n1936), .Q(n1934));
   XOR2X1 U1915 (.IN1(n1560), .IN2(n1561), .Q(n1110));
   XOR2X1 U1916 (.IN1(n1440), .IN2(n1138), .Q(n1561));
   XNOR2X1 U1917 (.IN1(n586), .IN2(n511), .Q(n1138));
   XNOR2X1 U1918 (.IN1(n518), .IN2(n572), .Q(n1560));
   XOR2X1 U1919 (.IN1(round_key[101]), .IN2(block[101]), .Q(n1929));
   AO221X1 U1920 (.IN1(n461), .IN2(new_sboxw[4]), .IN3(n664), .IN4(n1937), .IN5(n1938), .Q(
          n2128));
   OAI222X1 U1921 (.IN1(n1939), .IN2(n197), .IN3(n2218), .IN4(n1940), .IN5(n1941), .IN6(
          n926), .QN(n1938));
   XOR2X1 U1924 (.IN1(n548), .IN2(n562), .Q(n1124));
   XNOR2X1 U1925 (.IN1(n1348), .IN2(n1944), .Q(n562));
   XOR2X1 U1926 (.IN1(n1310), .IN2(n573), .Q(n548));
   XNOR2X1 U1927 (.IN1(n587), .IN2(n1288), .Q(n573));
   XNOR2X1 U1928 (.IN1(n1568), .IN2(n516), .Q(n531));
   XNOR2X1 U1929 (.IN1(n332), .IN2(round_key[99]), .Q(n578));
   XNOR2X1 U1930 (.IN1(n546), .IN2(n561), .Q(n1123));
   XNOR2X1 U1931 (.IN1(n1539), .IN2(n1945), .Q(n561));
   XOR2X1 U1932 (.IN1(n1537), .IN2(n1587), .Q(n546));
   XOR3X1 U1933 (.IN1(n555), .IN2(n540), .IN3(n1946), .Q(n1942));
   XOR2X1 U1934 (.IN1(n514), .IN2(n557), .Q(n1946));
   XOR2X1 U1935 (.IN1(n1136), .IN2(n618), .Q(n557));
   XNOR2X1 U1936 (.IN1(n302), .IN2(round_key[116]), .Q(n514));
   XNOR2X1 U1937 (.IN1(n1263), .IN2(new_block[124]), .Q(n540));
   XNOR2X1 U1938 (.IN1(n317), .IN2(round_key[108]), .Q(n555));
   XOR2X1 U1939 (.IN1(n1572), .IN2(n1573), .Q(n1120));
   XOR2X1 U1940 (.IN1(n539), .IN2(n1586), .Q(n1573));
   XOR2X1 U1941 (.IN1(n601), .IN2(n1093), .Q(n1586));
   XOR2X1 U1942 (.IN1(n1261), .IN2(n1584), .Q(n1572));
   XNOR2X1 U1943 (.IN1(n1161), .IN2(n518), .Q(n1584));
   XOR2X1 U1944 (.IN1(round_key[100]), .IN2(block[100]), .Q(n1937));
   AO221X1 U1945 (.IN1(n461), .IN2(new_sboxw[3]), .IN3(n679), .IN4(n1947), .IN5(n1948), .Q(
          n2129));
   OAI222X1 U1946 (.IN1(n1949), .IN2(n199), .IN3(n2220), .IN4(n1950), .IN5(n1951), .IN6(
          n926), .QN(n1948));
   XOR2X1 U1949 (.IN1(n579), .IN2(n1944), .Q(n1135));
   XNOR2X1 U1950 (.IN1(n602), .IN2(n1310), .Q(n1944));
   XOR2X1 U1951 (.IN1(n1348), .IN2(n605), .Q(n579));
   XNOR2X1 U1952 (.IN1(n592), .IN2(n516), .Q(n1587));
   XOR2X1 U1953 (.IN1(n333), .IN2(n1579), .Q(n592));
   XNOR2X1 U1954 (.IN1(n577), .IN2(n1945), .Q(n1134));
   XNOR2X1 U1955 (.IN1(n609), .IN2(n1537), .Q(n1945));
   XOR2X1 U1956 (.IN1(n1539), .IN2(n1604), .Q(n577));
   XOR3X1 U1957 (.IN1(n569), .IN2(n1136), .IN3(n1954), .Q(n1952));
   XOR2X1 U1958 (.IN1(n570), .IN2(n572), .Q(n1954));
   XOR2X1 U1959 (.IN1(n1149), .IN2(n618), .Q(n572));
   XOR2X1 U1960 (.IN1(n303), .IN2(n1371), .Q(n570));
   XOR2X1 U1961 (.IN1(round_key[123]), .IN2(new_block[123]), .Q(n1136));
   XOR2X1 U1962 (.IN1(n318), .IN2(n1470), .Q(n569));
   XOR2X1 U1963 (.IN1(n1583), .IN2(n1585), .Q(n1131));
   XNOR2X1 U1965 (.IN1(n620), .IN2(n511), .Q(n1163));
   XOR2X1 U1966 (.IN1(n1955), .IN2(n604), .Q(n1583));
   XOR2X1 U1967 (.IN1(round_key[99]), .IN2(block[99]), .Q(n1947));
   AO221X1 U1968 (.IN1(n461), .IN2(new_sboxw[2]), .IN3(n664), .IN4(n1956), .IN5(n1957), .Q(
          n2130));
   OAI222X1 U1969 (.IN1(n1958), .IN2(n200), .IN3(n2222), .IN4(n1959), .IN5(n1960), .IN6(
          n926), .QN(n1957));
   XNOR2X1 U1972 (.IN1(n605), .IN2(n594), .Q(n1148));
   XOR2X1 U1973 (.IN1(n621), .IN2(n508), .Q(n605));
   XNOR2X1 U1974 (.IN1(n1604), .IN2(n593), .Q(n1147));
   XOR2X1 U1975 (.IN1(n334), .IN2(n1594), .Q(n609));
   XOR3X1 U1976 (.IN1(n1149), .IN2(n586), .IN3(n1963), .Q(n1961));
   XOR2X1 U1977 (.IN1(n587), .IN2(n1161), .Q(n1963));
   XOR2X1 U1978 (.IN1(n304), .IN2(n1372), .Q(n587));
   XOR2X1 U1979 (.IN1(n319), .IN2(n1477), .Q(n586));
   XOR2X1 U1980 (.IN1(round_key[122]), .IN2(new_block[122]), .Q(n1149));
   XOR2X1 U1981 (.IN1(n1597), .IN2(n1598), .Q(n1144));
   XOR2X1 U1982 (.IN1(n1093), .IN2(n511), .Q(n1598));
   XOR2X1 U1983 (.IN1(new_block[111]), .IN2(round_key[111]), .Q(n511));
   XOR2X1 U1984 (.IN1(n1247), .IN2(n618), .Q(n1597));
   XOR2X1 U1985 (.IN1(round_key[98]), .IN2(block[98]), .Q(n1956));
   AO221X1 U1986 (.IN1(n461), .IN2(new_sboxw[1]), .IN3(n664), .IN4(n1964), .IN5(n1965), .Q(
          n2131));
   OAI222X1 U1987 (.IN1(n1966), .IN2(n201), .IN3(n2223), .IN4(n1967), .IN5(n1968), .IN6(
          n926), .QN(n1965));
   XOR2X1 U1990 (.IN1(n611), .IN2(n594), .Q(n1160));
   XOR2X1 U1991 (.IN1(n1310), .IN2(n1288), .Q(n594));
   XNOR2X1 U1992 (.IN1(n296), .IN2(round_key[119]), .Q(n508));
   XOR2X1 U1993 (.IN1(n610), .IN2(n593), .Q(n1159));
   XOR2X1 U1994 (.IN1(n1541), .IN2(n516), .Q(n593));
   XNOR2X1 U1995 (.IN1(n624), .IN2(n516), .Q(n1604));
   XOR2X1 U1996 (.IN1(n335), .IN2(n1595), .Q(n624));
   XOR3X1 U1997 (.IN1(n1161), .IN2(n601), .IN3(n1971), .Q(n1969));
   XNOR2X1 U1998 (.IN1(n602), .IN2(n604), .Q(n1971));
   XNOR2X1 U1999 (.IN1(n1173), .IN2(n618), .Q(n604));
   XOR2X1 U2000 (.IN1(n305), .IN2(n1377), .Q(n602));
   XNOR2X1 U2001 (.IN1(n321), .IN2(round_key[105]), .Q(n601));
   XOR2X1 U2002 (.IN1(round_key[121]), .IN2(new_block[121]), .Q(n1161));
   XOR2X1 U2003 (.IN1(n622), .IN2(n1616), .Q(n1156));
   XNOR2X1 U2004 (.IN1(n1440), .IN2(n539), .Q(n1616));
   XNOR2X1 U2005 (.IN1(n313), .IN2(round_key[110]), .Q(n1093));
   XOR2X1 U2006 (.IN1(n518), .IN2(n1955), .Q(n622));
   XOR2X1 U2007 (.IN1(n1248), .IN2(new_block[126]), .Q(n518));
   XOR2X1 U2008 (.IN1(round_key[97]), .IN2(block[97]), .Q(n1964));
   AO221X1 U2009 (.IN1(n461), .IN2(new_sboxw[0]), .IN3(n679), .IN4(n1972), .IN5(n1973), .Q(
          n2132));
   OAI222X1 U2010 (.IN1(n1974), .IN2(n202), .IN3(n2224), .IN4(n1975), .IN5(n1976), .IN6(
          n926), .QN(n1973));
   XOR3X1 U2012 (.IN1(n516), .IN2(n610), .IN3(n611), .Q(n1979));
   XNOR2X1 U2013 (.IN1(n509), .IN2(n542), .Q(n611));
   XNOR2X1 U2014 (.IN1(n300), .IN2(round_key[117]), .Q(n542));
   XNOR2X1 U2015 (.IN1(n298), .IN2(round_key[118]), .Q(n509));
   XNOR2X1 U2016 (.IN1(n1537), .IN2(n547), .Q(n610));
   XNOR2X1 U2017 (.IN1(n328), .IN2(round_key[101]), .Q(n547));
   XNOR2X1 U2018 (.IN1(n326), .IN2(round_key[102]), .Q(n1541));
   XOR2X1 U2019 (.IN1(new_block[103]), .IN2(round_key[103]), .Q(n516));
   XOR3X1 U2020 (.IN1(n618), .IN2(n1173), .IN3(n1936), .Q(n1978));
   XOR2X1 U2021 (.IN1(n539), .IN2(n1261), .Q(n1936));
   XOR2X1 U2022 (.IN1(n1262), .IN2(new_block[125]), .Q(n1955));
   XNOR2X1 U2023 (.IN1(n315), .IN2(round_key[109]), .Q(n539));
   XOR2X1 U2024 (.IN1(round_key[120]), .IN2(new_block[120]), .Q(n1173));
   XNOR2X1 U2025 (.IN1(n1231), .IN2(new_block[127]), .Q(n618));
   XOR2X1 U2027 (.IN1(n306), .IN2(n1382), .Q(n621));
   XOR2X1 U2028 (.IN1(n322), .IN2(n1520), .Q(n620));
   XOR2X1 U2029 (.IN1(round_key[96]), .IN2(block[96]), .Q(n1972));
   AO221X1 U2031 (.IN1(new_sboxw[0]), .IN2(n1088), .IN3(n785), .IN4(n1981), .IN5(n1982), .
          Q(n2133));
   OAI222X1 U2032 (.IN1(n1983), .IN2(n335), .IN3(n1595), .IN4(n1984), .IN5(n1985), .IN6(
          n926), .QN(n1982));
   XNOR2X1 U2035 (.IN1(n1870), .IN2(n905), .Q(n1067));
   XNOR2X1 U2036 (.IN1(n286), .IN2(round_key[69]), .Q(n905));
   XNOR2X1 U2037 (.IN1(n284), .IN2(round_key[70]), .Q(n890));
   XOR2X1 U2038 (.IN1(n1693), .IN2(n1703), .Q(n1064));
   XNOR2X1 U2039 (.IN1(n258), .IN2(round_key[85]), .Q(n917));
   XNOR2X1 U2040 (.IN1(n256), .IN2(round_key[86]), .Q(n901));
   XNOR2X1 U2041 (.IN1(n280), .IN2(round_key[71]), .Q(n990));
   XOR3X1 U2042 (.IN1(n1011), .IN2(n1531), .IN3(n1989), .Q(n1987));
   XOR2X1 U2043 (.IN1(n888), .IN2(n1623), .Q(n1989));
   XOR2X1 U2044 (.IN1(n1632), .IN2(new_block[93]), .Q(n1001));
   XOR2X1 U2045 (.IN1(round_key[95]), .IN2(new_block[95]), .Q(n888));
   XOR2X1 U2046 (.IN1(round_key[88]), .IN2(new_block[88]), .Q(n1531));
   XNOR2X1 U2047 (.IN1(n272), .IN2(round_key[77]), .Q(n1011));
   XOR2X1 U2048 (.IN1(n1075), .IN2(n1077), .Q(n1986));
   XOR2X1 U2049 (.IN1(n264), .IN2(n1744), .Q(n1077));
   XOR2X1 U2050 (.IN1(n278), .IN2(n1842), .Q(n1075));
   XOR2X1 U2051 (.IN1(round_key[64]), .IN2(block[64]), .Q(n1981));
   AND3X1 U2054 (.IN1(n520), .IN2(n436), .IN3(n926), .Q(n1375));
   AO21X1 U2056 (.IN1(ready), .IN2(n1994), .IN3(n833), .Q(n2134));
   AO221X1 U2057 (.IN1(n1992), .IN2(n2139), .IN3(round[3]), .IN4(n1996), .IN5(n2230), .Q(
          n2135));
   OR2X1 U2058 (.IN1(n1997), .IN2(round[2]), .Q(n1996));
   AO222X1 U2059 (.IN1(keylen), .IN2(n2230), .IN3(n1998), .IN4(n1999), .IN5(round[2]), .
          IN6(n1997), .Q(n2136));
   AO21X1 U2060 (.IN1(round[1]), .IN2(n2225), .IN3(n2000), .Q(n1997));
   AO221X1 U2061 (.IN1(n1999), .IN2(n203), .IN3(round[1]), .IN4(n2000), .IN5(n2230), .Q(
          n2137));
   AO21X1 U2062 (.IN1(round[0]), .IN2(n2225), .IN3(n2226), .Q(n2000));
   AO21X1 U2063 (.IN1(n2226), .IN2(round[0]), .IN3(n1999), .Q(n2138));
   AO21X1 U2065 (.IN1(n2002), .IN2(dec_ctrl_reg[1]), .IN3(n2227), .Q(n2140));
   AO22X1 U2067 (.IN1(n2004), .IN2(sword_ctr_reg[1]), .IN3(n2229), .IN4(n2005), .Q(n2141)
          );
   OR2X1 U2068 (.IN1(n1695), .IN2(n1376), .Q(n2005));
   AO22X1 U2069 (.IN1(n2004), .IN2(sword_ctr_reg[0]), .IN3(n2229), .IN4(n205), .Q(n2142)
          );
   AND2X1 U2070 (.IN1(n2002), .IN2(n1993), .Q(n2004));
   AND2X1 U2071 (.IN1(n2228), .IN2(n2003), .Q(n2002));
   aes_inv_sbox inv_sbox_inst (.sboxw(tmp_sboxw), .new_sboxw(new_sboxw));
   SDFFARX1 \block_w2_reg_reg[13]  (.D(n2087), .SI(new_block[44]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[45]), .QN(n227));
   SDFFARX1 \block_w2_reg_reg[12]  (.D(n2088), .SI(new_block[43]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[44]), .QN(n229));
   SDFFARX1 \block_w2_reg_reg[14]  (.D(n2086), .SI(new_block[45]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[46]), .QN(n225));
   SDFFARX1 \block_w0_reg_reg[19]  (.D(n2018), .SI(new_block[114]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[115]), .QN(n303));
   SDFFARX1 \block_w0_reg_reg[11]  (.D(n2026), .SI(new_block[106]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[107]), .QN(n318));
   SDFFARX1 \block_w1_reg_reg[12]  (.D(n2056), .SI(new_block[75]), .SE(test_se), .CLK(clk)
          , .RSTB(n1100), .Q(new_block[76]), .QN(n274));
   SDFFARX1 \block_w0_reg_reg[12]  (.D(n2025), .SI(new_block[107]), .SE(test_se), .CLK(clk)
          , .RSTB(n1180), .Q(new_block[108]), .QN(n317));
   SDFFARX1 \block_w0_reg_reg[22]  (.D(n2015), .SI(new_block[117]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[118]), .QN(n298));
   SDFFARX1 \block_w0_reg_reg[14]  (.D(n2023), .SI(new_block[109]), .SE(test_se), .CLK(clk)
          , .RSTB(n1192), .Q(new_block[110]), .QN(n313));
   SDFFARX1 \block_w0_reg_reg[4]  (.D(n2033), .SI(new_block[99]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[100]), .QN(n330));
   SDFFARX1 \block_w2_reg_reg[20]  (.D(n2080), .SI(new_block[51]), .SE(test_se), .CLK(clk)
          , .RSTB(n1133), .Q(new_block[52]), .QN(n215));
   SDFFARX1 \block_w2_reg_reg[4]  (.D(n2096), .SI(new_block[35]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[36]), .QN(n241));
   SDFFARX1 \block_w0_reg_reg[20]  (.D(n2017), .SI(new_block[115]), .SE(test_se), .CLK(clk)
          , .RSTB(n1112), .Q(new_block[116]), .QN(n302));
   SDFFARX1 \block_w2_reg_reg[5]  (.D(n2095), .SI(new_block[36]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[37]), .QN(n239));
   SDFFARX1 \block_w0_reg_reg[21]  (.D(n2016), .SI(new_block[116]), .SE(test_se), .CLK(clk)
          , .RSTB(n1125), .Q(new_block[117]), .QN(n300));
   SDFFARX1 \block_w1_reg_reg[13]  (.D(n2055), .SI(new_block[76]), .SE(test_se), .CLK(clk)
          , .RSTB(n1146), .Q(new_block[77]), .QN(n272));
   SDFFARX1 \block_w3_reg_reg[30]  (.D(n2102), .SI(n2238), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[30]), .QN(n2237));
   SDFFARX1 \block_w1_reg_reg[30]  (.D(n2038), .SI(n2254), .SE(test_se), .CLK(clk), .RSTB(
          n1192), .Q(new_block[94]), .QN(n2253));
   SDFFARX1 \block_w1_reg_reg[29]  (.D(n2039), .SI(n2255), .SE(test_se), .CLK(clk), .RSTB(
          n1125), .Q(new_block[93]), .QN(n2254));
   SDFFARX1 \block_w2_reg_reg[29]  (.D(n2071), .SI(n2247), .SE(test_se), .CLK(clk), .RSTB(
          n1169), .Q(new_block[61]), .QN(n2246));
   SDFFARX1 \block_w2_reg_reg[27]  (.D(n2073), .SI(n2249), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[59]), .QN(n2248));
   SDFFARX1 \block_w3_reg_reg[25]  (.D(n2107), .SI(n2243), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(new_block[25]), .QN(n2242));
   SDFFARX1 \block_w1_reg_reg[28]  (.D(n2040), .SI(n2256), .SE(test_se), .CLK(clk), .RSTB(
          n1133), .Q(new_block[92]), .QN(n2255));
   SDFFARX1 \block_w1_reg_reg[25]  (.D(n2043), .SI(n2259), .SE(test_se), .CLK(clk), .RSTB(
          n1203), .Q(new_block[89]), .QN(n2258));
   SDFFARX1 \block_w3_reg_reg[28]  (.D(n2104), .SI(n2240), .SE(test_se), .CLK(clk), .RSTB(
          n1099), .Q(new_block[28]), .QN(n2239));
   SDFFARX1 \block_w2_reg_reg[28]  (.D(n2072), .SI(n2248), .SE(test_se), .CLK(clk), .RSTB(
          n1180), .Q(new_block[60]), .QN(n2247));
   SDFFARX1 \block_w0_reg_reg[13]  (.D(n2024), .SI(new_block[108]), .SE(test_se), .CLK(clk)
          , .RSTB(n1169), .Q(new_block[109]), .QN(n315));
   SDFFARX1 \block_w3_reg_reg[29]  (.D(n2103), .SI(n2239), .SE(test_se), .CLK(clk), .RSTB(
          n1133), .Q(new_block[29]), .QN(n2238));
   SDFFARX1 \dec_ctrl_reg_reg[0]  (.D(n2139), .SI(n2236), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(dec_ctrl_reg[0]), .QN(n159));
   SDFFARX1 \dec_ctrl_reg_reg[1]  (.D(n2140), .SI(dec_ctrl_reg[0]), .SE(test_se), .CLK(clk)
          , .RSTB(n1089), .Q(dec_ctrl_reg[1]), .QN(n158));
   SDFFARX1 \round_ctr_reg_reg[0]  (.D(n2138), .SI(n2235), .SE(test_se), .CLK(clk), .RSTB(
          n1089), .Q(round[0]), .QN(n2234));
   NAND3X0 U140 (.IN1(n205), .IN2(n204), .IN3(n1374), .QN(n497));
   AND2X1 U141 (.IN1(n1375), .IN2(n496), .Q(n1));
   INVX0 U142 (.INP(n2), .ZN(n1087));
   NBUFFX2 U143 (.INP(n1076), .Z(n926));
   INVX0 U144 (.INP(n2), .ZN(n1081));
   INVX0 U145 (.INP(n2), .ZN(n1088));
   NBUFFX2 U146 (.INP(n1047), .Z(n1008));
   NBUFFX2 U147 (.INP(n1060), .Z(n985));
   NBUFFX2 U148 (.INP(n1060), .Z(n996));
   NBUFFX2 U149 (.INP(n1060), .Z(n979));
   NBUFFX2 U150 (.INP(n1047), .Z(n1022));
   NBUFFX2 U151 (.INP(n1047), .Z(n1033));
   NBUFFX2 U152 (.INP(n1076), .Z(n971));
   NBUFFX2 U153 (.INP(n1076), .Z(n939));
   NBUFFX2 U154 (.INP(n1205), .Z(n1193));
   NBUFFX2 U155 (.INP(n1205), .Z(n1192));
   NBUFFX2 U156 (.INP(n1216), .Z(n1146));
   NBUFFX2 U157 (.INP(n1217), .Z(n1125));
   NBUFFX2 U158 (.INP(n1217), .Z(n1112));
   NBUFFX2 U159 (.INP(n1218), .Z(n1100));
   NBUFFX2 U160 (.INP(n1216), .Z(n1180));
   NBUFFX2 U161 (.INP(n1216), .Z(n1169));
   NBUFFX2 U162 (.INP(n1218), .Z(n1099));
   NBUFFX2 U163 (.INP(n1217), .Z(n1133));
   NBUFFX2 U164 (.INP(n1218), .Z(n1089));
   NBUFFX2 U165 (.INP(n1205), .Z(n1203));
   XNOR2X1 U166 (.IN1(n1013), .IN2(n1025), .Q(n928));
   XNOR2X1 U167 (.IN1(n1207), .IN2(n1220), .Q(n681));
   XNOR2X1 U168 (.IN1(n1015), .IN2(n1027), .Q(n927));
   NAND2X0 U169 (.IN1(n1374), .IN2(n619), .QN(n2));
   NBUFFX2 U170 (.INP(n505), .Z(n1076));
   NAND2X1 U171 (.IN1(n1374), .IN2(n457), .QN(n3));
   INVX0 U172 (.INP(n498), .ZN(n456));
   NAND2X1 U173 (.IN1(n1374), .IN2(n538), .QN(n4));
   NAND2X1 U174 (.IN1(n1374), .IN2(n462), .QN(n142));
   NBUFFX2 U175 (.INP(n505), .Z(n1060));
   NBUFFX2 U176 (.INP(n505), .Z(n1047));
   NBUFFX2 U177 (.INP(reset_n), .Z(n1216));
   NBUFFX2 U178 (.INP(reset_n), .Z(n1205));
   NBUFFX2 U179 (.INP(reset_n), .Z(n1218));
   NBUFFX2 U180 (.INP(reset_n), .Z(n1217));
   INVX0 U181 (.INP(n1239), .ZN(n2199));
   INVX0 U182 (.INP(n1791), .ZN(n2156));
   XNOR2X1 U183 (.IN1(n1210), .IN2(n2181), .Q(n1209));
   INVX0 U184 (.INP(n1903), .ZN(n1771));
   XNOR2X1 U185 (.IN1(n1210), .IN2(n1224), .Q(n682));
   INVX0 U186 (.INP(n1278), .ZN(n2202));
   INVX0 U187 (.INP(n1195), .ZN(n2213));
   INVX0 U188 (.INP(n860), .ZN(n2155));
   INVX0 U189 (.INP(n1853), .ZN(n1764));
   INVX0 U190 (.INP(n1223), .ZN(n2200));
   INVX0 U191 (.INP(n1562), .ZN(n1399));
   XNOR2X1 U192 (.IN1(n1666), .IN2(n1731), .Q(n1233));
   XNOR2X1 U193 (.IN1(n1502), .IN2(n1874), .Q(n1037));
   INVX0 U194 (.INP(n1067), .ZN(n1863));
   INVX0 U195 (.INP(n1452), .ZN(n2158));
   INVX0 U196 (.INP(n1616), .ZN(n1416));
   INVX0 U197 (.INP(n772), .ZN(n2167));
   XNOR2X1 U198 (.IN1(n143), .IN2(n526), .Q(n524));
   XNOR3X1 U199 (.IN1(n529), .IN2(n1348), .IN3(n530), .Q(n143));
   INVX0 U200 (.INP(n1268), .ZN(n2198));
   INVX0 U201 (.INP(n903), .ZN(n1613));
   INVX0 U202 (.INP(n1163), .ZN(n1391));
   XNOR2X1 U203 (.IN1(n1480), .IN2(n1479), .Q(n912));
   INVX0 U204 (.INP(n1138), .ZN(n1392));
   INVX0 U205 (.INP(n1501), .ZN(n1760));
   INVX0 U206 (.INP(n929), .ZN(n1861));
   OR2X1 U207 (.IN1(n1990), .IN2(n1991), .Q(n505));
   INVX0 U208 (.INP(n2139), .ZN(n2226));
   AND2X1 U209 (.IN1(n1375), .IN2(n499), .Q(n144));
   INVX0 U210 (.INP(n2001), .ZN(n2225));
   INVX0 U211 (.INP(round_key[10]), .ZN(n2209));
   XNOR2X1 U212 (.IN1(n145), .IN2(n1720), .Q(n1718));
   XNOR3X1 U213 (.IN1(n1206), .IN2(n1210), .IN3(n1721), .Q(n145));
   XNOR2X1 U214 (.IN1(n146), .IN2(n1727), .Q(n1725));
   XNOR3X1 U215 (.IN1(n1219), .IN2(n1224), .IN3(n1729), .Q(n146));
   INVX0 U216 (.INP(round_key[42]), .ZN(n2163));
   XOR2X1 U217 (.IN1(n147), .IN2(n148), .Q(n784));
   XNOR3X1 U218 (.IN1(n791), .IN2(n792), .IN3(n793), .Q(n147));
   XNOR3X1 U219 (.IN1(n787), .IN2(n788), .IN3(n789), .Q(n148));
   XNOR2X1 U220 (.IN1(n1406), .IN2(n149), .Q(n1405));
   XNOR3X1 U221 (.IN1(n790), .IN2(n809), .IN3(n1408), .Q(n149));
   INVX0 U222 (.INP(round_key[23]), .ZN(n2189));
   XOR3X1 U223 (.IN1(n150), .IN2(n1204), .IN3(n151), .Q(n1202));
   XNOR3X1 U224 (.IN1(n633), .IN2(n649), .IN3(n1209), .Q(n150));
   XNOR3X1 U225 (.IN1(n1206), .IN2(n1207), .IN3(n1208), .Q(n151));
   INVX0 U226 (.INP(round_key[2]), .ZN(n2222));
   XNOR2X1 U227 (.IN1(n663), .IN2(n152), .Q(n662));
   XNOR3X1 U228 (.IN1(n665), .IN2(n2205), .IN3(n666), .Q(n152));
   XNOR2X1 U229 (.IN1(n1641), .IN2(n153), .Q(n1640));
   XNOR3X1 U230 (.IN1(n1643), .IN2(n2205), .IN3(n666), .Q(n153));
   INVX0 U231 (.INP(n899), .ZN(n1772));
   XNOR2X1 U232 (.IN1(n154), .IN2(n1061), .Q(n1059));
   XNOR3X1 U233 (.IN1(n1064), .IN2(n1065), .IN3(n1066), .Q(n154));
   XNOR2X1 U234 (.IN1(n1021), .IN2(n155), .Q(n1020));
   XNOR3X1 U235 (.IN1(n884), .IN2(n930), .IN3(n1023), .Q(n155));
   INVX0 U236 (.INP(round_key[22]), .ZN(n2190));
   XNOR3X1 U237 (.IN1(n678), .IN2(n156), .IN3(n680), .Q(n677));
   XNOR3X1 U238 (.IN1(n633), .IN2(n2183), .IN3(n683), .Q(n156));
   XNOR3X1 U239 (.IN1(n678), .IN2(n1650), .IN3(n157), .Q(n1649));
   XNOR3X1 U240 (.IN1(n681), .IN2(n1195), .IN3(n682), .Q(n157));
   INVX0 U241 (.INP(n901), .ZN(n1693));
   XNOR3X1 U242 (.IN1(n924), .IN2(n160), .IN3(n1487), .Q(n1485));
   XNOR3X1 U243 (.IN1(n884), .IN2(n1634), .IN3(n1488), .Q(n160));
   XNOR3X1 U244 (.IN1(n924), .IN2(n925), .IN3(n161), .Q(n923));
   XNOR3X1 U245 (.IN1(n927), .IN2(n1861), .IN3(n928), .Q(n161));
   INVX0 U246 (.INP(n655), .ZN(n2215));
   INVX0 U247 (.INP(n890), .ZN(n1870));
   XNOR2X1 U248 (.IN1(n790), .IN2(n806), .Q(n774));
   INVX0 U249 (.INP(round_key[43]), .ZN(n2162));
   XNOR3X1 U250 (.IN1(n751), .IN2(n767), .IN3(n162), .Q(n766));
   XNOR2X1 U251 (.IN1(n769), .IN2(n770), .Q(n162));
   INVX0 U252 (.INP(n648), .ZN(n2203));
   XNOR2X1 U253 (.IN1(n163), .IN2(n1753), .Q(n1751));
   XNOR3X1 U254 (.IN1(n739), .IN2(n1264), .IN3(n1755), .Q(n163));
   INVX0 U255 (.INP(n1236), .ZN(n2221));
   XNOR2X1 U256 (.IN1(n165), .IN2(n647), .Q(n645));
   XNOR3X1 U257 (.IN1(n652), .IN2(n653), .IN3(n654), .Q(n165));
   INVX0 U258 (.INP(round_key[17]), .ZN(n2195));
   INVX0 U259 (.INP(round_key[18]), .ZN(n2194));
   XNOR3X1 U260 (.IN1(n799), .IN2(n168), .IN3(n801), .Q(n798));
   XNOR2X1 U261 (.IN1(n755), .IN2(n2167), .Q(n168));
   XNOR2X1 U262 (.IN1(n771), .IN2(n2155), .Q(n1423));
   INVX0 U263 (.INP(round_key[40]), .ZN(n2165));
   XNOR2X1 U264 (.IN1(n174), .IN2(n1417), .Q(n1415));
   XNOR3X1 U265 (.IN1(n818), .IN2(n819), .IN3(n1420), .Q(n174));
   XNOR2X1 U266 (.IN1(n1398), .IN2(n175), .Q(n1397));
   XNOR3X1 U267 (.IN1(n1400), .IN2(n2149), .IN3(n789), .Q(n175));
   XNOR3X1 U268 (.IN1(n176), .IN2(n178), .IN3(n179), .Q(n1215));
   XNOR3X1 U269 (.IN1(n1222), .IN2(n1223), .IN3(n1224), .Q(n176));
   XNOR2X1 U270 (.IN1(n1184), .IN2(n2213), .Q(n178));
   XNOR3X1 U271 (.IN1(n1219), .IN2(n1220), .IN3(n1221), .Q(n179));
   INVX0 U272 (.INP(round_key[74]), .ZN(n1826));
   XNOR2X1 U273 (.IN1(n181), .IN2(n1009), .Q(n1007));
   XNOR3X1 U274 (.IN1(n1012), .IN2(n1013), .IN3(n1014), .Q(n181));
   INVX0 U275 (.INP(round_key[75]), .ZN(n1817));
   XNOR2X1 U276 (.IN1(n183), .IN2(n997), .Q(n995));
   XNOR3X1 U277 (.IN1(n1000), .IN2(n1001), .IN3(n1002), .Q(n183));
   INVX0 U278 (.INP(round_key[11]), .ZN(n2208));
   XNOR2X1 U279 (.IN1(n189), .IN2(n1710), .Q(n1708));
   XNOR3X1 U280 (.IN1(n1194), .IN2(n1712), .IN3(n1713), .Q(n189));
   XNOR3X1 U281 (.IN1(n815), .IN2(n191), .IN3(n817), .Q(n814));
   XNOR2X1 U282 (.IN1(n821), .IN2(n822), .Q(n191));
   XNOR3X1 U283 (.IN1(n695), .IN2(n696), .IN3(n192), .Q(n691));
   XNOR2X1 U284 (.IN1(n2199), .IN2(n698), .Q(n192));
   INVX0 U285 (.INP(round_key[73]), .ZN(n1834));
   XNOR2X1 U286 (.IN1(n555), .IN2(n1399), .Q(n528));
   INVX0 U287 (.INP(round_key[107]), .ZN(n1470));
   XOR2X1 U288 (.IN1(n194), .IN2(n196), .Q(n1547));
   XNOR3X1 U289 (.IN1(n532), .IN2(n547), .IN3(n529), .Q(n194));
   XNOR3X1 U290 (.IN1(n1550), .IN2(n518), .IN3(n528), .Q(n196));
   INVX0 U291 (.INP(n756), .ZN(n2143));
   INVX0 U292 (.INP(round_key[9]), .ZN(n2210));
   INVX0 U293 (.INP(round_key[81]), .ZN(n1738));
   INVX0 U294 (.INP(round_key[65]), .ZN(n1902));
   INVX0 U295 (.INP(round_key[1]), .ZN(n2223));
   INVX0 U296 (.INP(round_key[106]), .ZN(n1477));
   XNOR3X1 U297 (.IN1(n517), .IN2(n531), .IN3(n198), .Q(n1567));
   XNOR2X1 U298 (.IN1(n1569), .IN2(n1570), .Q(n198));
   XNOR3X1 U299 (.IN1(n517), .IN2(n547), .IN3(n206), .Q(n1555));
   XNOR2X1 U300 (.IN1(n1557), .IN2(n1558), .Q(n206));
   INVX0 U301 (.INP(n917), .ZN(n1703));
   INVX0 U302 (.INP(n905), .ZN(n1872));
   INVX0 U303 (.INP(n671), .ZN(n2217));
   INVX0 U304 (.INP(n758), .ZN(n2159));
   XNOR3X1 U305 (.IN1(n695), .IN2(n1241), .IN3(n207), .Q(n1737));
   XNOR2X1 U306 (.IN1(n1665), .IN2(n698), .Q(n207));
   XNOR2X1 U307 (.IN1(n208), .IN2(n1034), .Q(n1032));
   XNOR3X1 U308 (.IN1(n1037), .IN2(n1038), .IN3(n1039), .Q(n208));
   XNOR3X1 U309 (.IN1(n690), .IN2(n1660), .IN3(n210), .Q(n1659));
   XOR3X1 U310 (.IN1(n693), .IN2(n1237), .IN3(n694), .Q(n210));
   INVX0 U311 (.INP(n1541), .ZN(n1537));
   INVX0 U312 (.INP(n651), .ZN(n2205));
   INVX0 U313 (.INP(round_key[8]), .ZN(n2211));
   INVX0 U314 (.INP(n1875), .ZN(n1614));
   XNOR2X1 U315 (.IN1(n212), .IN2(n1048), .Q(n1046));
   XNOR3X1 U316 (.IN1(n1050), .IN2(n1051), .IN3(n1052), .Q(n212));
   INVX0 U317 (.INP(round_key[94]), .ZN(n1615));
   XNOR3X1 U318 (.IN1(n1230), .IN2(n214), .IN3(n1232), .Q(n1229));
   XNOR2X1 U319 (.IN1(n1236), .IN2(n1237), .Q(n214));
   XNOR3X1 U320 (.IN1(n1882), .IN2(n220), .IN3(n1884), .Q(n1881));
   XNOR2X1 U321 (.IN1(n1041), .IN2(n941), .Q(n220));
   XNOR3X1 U322 (.IN1(n969), .IN2(n1519), .IN3(n221), .Q(n1518));
   XNOR3X1 U323 (.IN1(n956), .IN2(n973), .IN3(n974), .Q(n221));
   XNOR3X1 U324 (.IN1(n969), .IN2(n970), .IN3(n223), .Q(n968));
   XNOR3X1 U325 (.IN1(n972), .IN2(n973), .IN3(n974), .Q(n223));
   INVX0 U326 (.INP(n1712), .ZN(n2181));
   INVX0 U327 (.INP(round_key[29]), .ZN(n2182));
   INVX0 U328 (.INP(round_key[64]), .ZN(n1910));
   XNOR3X1 U329 (.IN1(n937), .IN2(n1496), .IN3(n224), .Q(n1495));
   XOR3X1 U330 (.IN1(n940), .IN2(n1041), .IN3(n942), .Q(n224));
   XNOR3X1 U331 (.IN1(n937), .IN2(n938), .IN3(n226), .Q(n936));
   XOR3X1 U332 (.IN1(n940), .IN2(n941), .IN3(n942), .Q(n226));
   INVX0 U333 (.INP(round_key[0]), .ZN(n2224));
   INVX0 U334 (.INP(n775), .ZN(n2145));
   XNOR3X1 U335 (.IN1(n790), .IN2(n808), .IN3(n228), .Q(n1797));
   XNOR2X1 U336 (.IN1(n806), .IN2(n776), .Q(n228));
   XNOR3X1 U337 (.IN1(n1322), .IN2(n1323), .IN3(n235), .Q(n1321));
   XNOR3X1 U338 (.IN1(n1325), .IN2(n772), .IN3(n1326), .Q(n235));
   INVX0 U339 (.INP(round_key[82]), .ZN(n1726));
   XNOR3X1 U340 (.IN1(n912), .IN2(n236), .IN3(n1478), .Q(n1476));
   XNOR3X1 U341 (.IN1(n884), .IN2(n930), .IN3(n918), .Q(n236));
   XNOR3X1 U342 (.IN1(n912), .IN2(n913), .IN3(n238), .Q(n911));
   XNOR3X1 U343 (.IN1(n915), .IN2(n1892), .IN3(n916), .Q(n238));
   XNOR3X1 U344 (.IN1(n1120), .IN2(n1942), .IN3(n240), .Q(n1941));
   XOR3X1 U345 (.IN1(n1123), .IN2(n531), .IN3(n1124), .Q(n240));
   XNOR3X1 U346 (.IN1(n242), .IN2(n247), .IN3(n248), .Q(n1899));
   XNOR3X1 U347 (.IN1(n963), .IN2(n977), .IN3(n1904), .Q(n242));
   XNOR2X1 U348 (.IN1(n956), .IN2(n972), .Q(n247));
   XNOR3X1 U349 (.IN1(n1067), .IN2(n1065), .IN3(n1068), .Q(n248));
   XNOR3X1 U350 (.IN1(n1891), .IN2(n249), .IN3(n1893), .Q(n1890));
   XNOR2X1 U351 (.IN1(n1053), .IN2(n956), .Q(n249));
   INVX0 U352 (.INP(round_key[66]), .ZN(n1901));
   XNOR3X1 U353 (.IN1(n250), .IN2(n1789), .IN3(n1790), .Q(n1787));
   XNOR2X1 U354 (.IN1(n1315), .IN2(n1316), .Q(n250));
   XNOR3X1 U355 (.IN1(n1309), .IN2(n251), .IN3(n1311), .Q(n1308));
   XNOR3X1 U356 (.IN1(n1314), .IN2(n808), .IN3(n1315), .Q(n251));
   INVX0 U357 (.INP(round_key[34]), .ZN(n2176));
   INVX0 U358 (.INP(round_key[48]), .ZN(n2153));
   XNOR3X1 U359 (.IN1(n1338), .IN2(n825), .IN3(n252), .Q(n1807));
   XNOR2X1 U360 (.IN1(n1791), .IN2(n1419), .Q(n252));
   INVX0 U361 (.INP(round_key[16]), .ZN(n2196));
   INVX0 U362 (.INP(round_key[72]), .ZN(n1842));
   XNOR2X1 U363 (.IN1(n539), .IN2(n1163), .Q(n1585));
   INVX0 U364 (.INP(round_key[104]), .ZN(n1520));
   XOR3X1 U365 (.IN1(n578), .IN2(n1587), .IN3(n254), .Q(n1578));
   XNOR2X1 U366 (.IN1(n1580), .IN2(n1581), .Q(n254));
   XNOR3X1 U367 (.IN1(n555), .IN2(n540), .IN3(n255), .Q(n1121));
   XNOR2X1 U368 (.IN1(n1399), .IN2(n532), .Q(n255));
   INVX0 U369 (.INP(n751), .ZN(n2169));
   XNOR3X1 U370 (.IN1(n257), .IN2(n259), .IN3(n266), .Q(n1869));
   XNOR3X1 U371 (.IN1(n1876), .IN2(n1853), .IN3(n1025), .Q(n257));
   XNOR2X1 U372 (.IN1(n989), .IN2(n929), .Q(n259));
   XNOR3X1 U373 (.IN1(n1024), .IN2(n1027), .IN3(n1028), .Q(n266));
   INVX0 U374 (.INP(round_key[67]), .ZN(n1900));
   XNOR3X1 U375 (.IN1(n917), .IN2(n1614), .IN3(n267), .Q(n1469));
   XNOR2X1 U376 (.IN1(n899), .IN2(n1764), .Q(n267));
   XNOR2X1 U377 (.IN1(n268), .IN2(n898), .Q(n896));
   XNOR3X1 U378 (.IN1(n902), .IN2(n903), .IN3(n904), .Q(n268));
   XNOR2X1 U379 (.IN1(n1439), .IN2(n269), .Q(n1438));
   XNOR3X1 U380 (.IN1(n843), .IN2(n858), .IN3(n1441), .Q(n269));
   INVX0 U381 (.INP(n1810), .ZN(n1926));
   INVX0 U382 (.INP(round_key[61]), .ZN(n1935));
   INVX0 U383 (.INP(n1093), .ZN(n1440));
   XNOR2X1 U384 (.IN1(n271), .IN2(n1607), .Q(n1605));
   XNOR3X1 U385 (.IN1(n611), .IN2(n610), .IN3(n607), .Q(n271));
   INVX0 U386 (.INP(n777), .ZN(n1912));
   INVX0 U387 (.INP(round_key[62]), .ZN(n1919));
   INVX0 U388 (.INP(n767), .ZN(n2171));
   XNOR3X1 U389 (.IN1(n1358), .IN2(n1359), .IN3(n273), .Q(n1357));
   XOR3X1 U390 (.IN1(n856), .IN2(n1361), .IN3(n1362), .Q(n273));
   XNOR3X1 U391 (.IN1(n857), .IN2(n843), .IN3(n279), .Q(n1824));
   XNOR2X1 U392 (.IN1(n860), .IN2(n1442), .Q(n279));
   XNOR2X1 U393 (.IN1(n281), .IN2(n554), .Q(n552));
   XOR3X1 U394 (.IN1(n558), .IN2(n559), .IN3(n560), .Q(n281));
   XNOR3X1 U395 (.IN1(n282), .IN2(n283), .IN3(n285), .Q(n1260));
   XNOR3X1 U396 (.IN1(n726), .IN2(n714), .IN3(n1267), .Q(n282));
   XNOR2X1 U397 (.IN1(n723), .IN2(n1266), .Q(n283));
   XNOR3X1 U398 (.IN1(n738), .IN2(n1264), .IN3(n1265), .Q(n285));
   INVX0 U399 (.INP(n508), .ZN(n1288));
   XNOR3X1 U400 (.IN1(n1110), .IN2(n1111), .IN3(n287), .Q(n1109));
   XNOR3X1 U401 (.IN1(n1113), .IN2(n1539), .IN3(n1114), .Q(n287));
   XNOR3X1 U402 (.IN1(n1110), .IN2(n1934), .IN3(n293), .Q(n1933));
   XNOR3X1 U403 (.IN1(n1113), .IN2(n1549), .IN3(n1114), .Q(n293));
   XNOR3X1 U404 (.IN1(n294), .IN2(n851), .IN3(n852), .Q(n849));
   XNOR3X1 U405 (.IN1(n857), .IN2(n858), .IN3(n859), .Q(n294));
   XNOR3X1 U406 (.IN1(n720), .IN2(n295), .IN3(n1683), .Q(n1681));
   XNOR3X1 U407 (.IN1(n726), .IN2(n713), .IN3(n1684), .Q(n295));
   XNOR3X1 U408 (.IN1(n726), .IN2(n713), .IN3(n297), .Q(n721));
   XNOR2X1 U409 (.IN1(n2198), .IN2(n728), .Q(n297));
   XNOR3X1 U410 (.IN1(n299), .IN2(n301), .IN3(n308), .Q(n831));
   XNOR3X1 U411 (.IN1(n840), .IN2(n841), .IN3(n842), .Q(n299));
   XNOR2X1 U412 (.IN1(n838), .IN2(n839), .Q(n301));
   XOR3X1 U413 (.IN1(n835), .IN2(n836), .IN3(n837), .Q(n308));
   XOR3X1 U414 (.IN1(n309), .IN2(n1633), .IN3(n310), .Q(n1631));
   XNOR2X1 U415 (.IN1(n652), .IN2(n656), .Q(n309));
   XNOR3X1 U416 (.IN1(n671), .IN2(n2181), .IN3(n657), .Q(n310));
   INVX0 U417 (.INP(n1001), .ZN(n1623));
   INVX0 U418 (.INP(round_key[93]), .ZN(n1632));
   XNOR3X1 U419 (.IN1(n756), .IN2(n760), .IN3(n311), .Q(n1449));
   XNOR2X1 U420 (.IN1(n791), .IN2(n1373), .Q(n311));
   INVX0 U421 (.INP(n821), .ZN(n2175));
   XNOR3X1 U422 (.IN1(n312), .IN2(n1780), .IN3(n1781), .Q(n1778));
   XNOR2X1 U423 (.IN1(n1912), .IN2(n791), .Q(n312));
   XNOR3X1 U424 (.IN1(n314), .IN2(n1298), .IN3(n1299), .Q(n1296));
   XNOR2X1 U425 (.IN1(n1303), .IN2(n1912), .Q(n314));
   INVX0 U426 (.INP(round_key[80]), .ZN(n1744));
   INVX0 U427 (.INP(round_key[21]), .ZN(n2191));
   INVX0 U428 (.INP(round_key[32]), .ZN(n2178));
   INVX0 U429 (.INP(round_key[98]), .ZN(n1579));
   INVX0 U430 (.INP(round_key[96]), .ZN(n1595));
   INVX0 U431 (.INP(n1011), .ZN(n1788));
   XNOR2X1 U432 (.IN1(n537), .IN2(n316), .Q(n536));
   XNOR3X1 U433 (.IN1(n539), .IN2(n540), .IN3(n541), .Q(n316));
   XNOR2X1 U434 (.IN1(n320), .IN2(n754), .Q(n752));
   XNOR3X1 U435 (.IN1(n2149), .IN2(n760), .IN3(n761), .Q(n320));
   INVX0 U436 (.INP(round_key[97]), .ZN(n1594));
   INVX0 U437 (.INP(round_key[41]), .ZN(n2164));
   INVX0 U438 (.INP(round_key[50]), .ZN(n2151));
   INVX0 U439 (.INP(n518), .ZN(n1247));
   XOR2X1 U440 (.IN1(n324), .IN2(n325), .Q(n1593));
   XOR3X1 U441 (.IN1(n594), .IN2(n593), .IN3(n590), .Q(n324));
   XNOR3X1 U442 (.IN1(n1596), .IN2(n1497), .IN3(n589), .Q(n325));
   INVX0 U443 (.INP(round_key[126]), .ZN(n1248));
   XNOR3X1 U444 (.IN1(n888), .IN2(n1075), .IN3(n327), .Q(n1074));
   XNOR2X1 U445 (.IN1(n886), .IN2(n917), .Q(n327));
   INVX0 U446 (.INP(n1955), .ZN(n1261));
   INVX0 U447 (.INP(round_key[125]), .ZN(n1262));
   INVX0 U448 (.INP(round_key[30]), .ZN(n2180));
   INVX0 U449 (.INP(n547), .ZN(n1539));
   XNOR3X1 U450 (.IN1(n329), .IN2(n331), .IN3(n336), .Q(n1860));
   XNOR3X1 U451 (.IN1(n1864), .IN2(n1001), .IN3(n1013), .Q(n329));
   XNOR2X1 U452 (.IN1(n905), .IN2(n989), .Q(n331));
   XNOR3X1 U453 (.IN1(n1012), .IN2(n1015), .IN3(n1016), .Q(n336));
   INVX0 U454 (.INP(n791), .ZN(n2147));
   XOR3X1 U455 (.IN1(n337), .IN2(n338), .IN3(n1101), .Q(n1098));
   XNOR2X1 U456 (.IN1(n557), .IN2(n542), .Q(n337));
   XNOR3X1 U457 (.IN1(n539), .IN2(n1247), .IN3(n1104), .Q(n338));
   XOR2X1 U458 (.IN1(n667), .IN2(n684), .Q(n652));
   INVX0 U459 (.INP(round_key[49]), .ZN(n2152));
   XNOR3X1 U460 (.IN1(n1850), .IN2(n1851), .IN3(n339), .Q(n1849));
   XNOR3X1 U461 (.IN1(n1000), .IN2(n1788), .IN3(n1003), .Q(n339));
   XNOR2X1 U462 (.IN1(n340), .IN2(n1761), .Q(n1759));
   XOR3X1 U463 (.IN1(n1279), .IN2(n1277), .IN3(n1763), .Q(n340));
   XOR3X1 U464 (.IN1(n1191), .IN2(n341), .IN3(n342), .Q(n1190));
   XNOR2X1 U465 (.IN1(n671), .IN2(n655), .Q(n341));
   XNOR3X1 U466 (.IN1(n1194), .IN2(n1195), .IN3(n1196), .Q(n342));
   XNOR2X1 U467 (.IN1(n343), .IN2(n568), .Q(n566));
   XNOR3X1 U468 (.IN1(n574), .IN2(n575), .IN3(n576), .Q(n343));
   INVX0 U469 (.INP(round_key[33]), .ZN(n2177));
   XNOR3X1 U470 (.IN1(n1131), .IN2(n1132), .IN3(n344), .Q(n1130));
   XNOR3X1 U471 (.IN1(n1134), .IN2(n1568), .IN3(n1135), .Q(n344));
   INVX0 U472 (.INP(round_key[112]), .ZN(n1382));
   XNOR3X1 U473 (.IN1(n1131), .IN2(n1952), .IN3(n345), .Q(n1951));
   XNOR3X1 U474 (.IN1(n1134), .IN2(n1587), .IN3(n1135), .Q(n345));
   XNOR2X1 U475 (.IN1(n346), .IN2(n1745), .Q(n1743));
   XNOR3X1 U476 (.IN1(n1255), .IN2(n1251), .IN3(n1747), .Q(n346));
   XNOR2X1 U477 (.IN1(n347), .IN2(n600), .Q(n598));
   XOR3X1 U478 (.IN1(n606), .IN2(n607), .IN3(n608), .Q(n347));
   XNOR3X1 U479 (.IN1(n704), .IN2(n705), .IN3(n348), .Q(n703));
   XNOR3X1 U480 (.IN1(n707), .IN2(n708), .IN3(n709), .Q(n348));
   XNOR3X1 U481 (.IN1(n704), .IN2(n1673), .IN3(n349), .Q(n1672));
   XNOR3X1 U482 (.IN1(n723), .IN2(n708), .IN3(n709), .Q(n349));
   INVX0 U483 (.INP(n509), .ZN(n1310));
   XNOR3X1 U484 (.IN1(n1156), .IN2(n1969), .IN3(n350), .Q(n1968));
   XOR3X1 U485 (.IN1(n1604), .IN2(n1159), .IN3(n1160), .Q(n350));
   XOR3X1 U486 (.IN1(n351), .IN2(n352), .IN3(n1249), .Q(n1246));
   XNOR3X1 U487 (.IN1(n711), .IN2(n1253), .IN3(n1254), .Q(n351));
   XNOR2X1 U488 (.IN1(n707), .IN2(n723), .Q(n352));
   XNOR3X1 U489 (.IN1(n1346), .IN2(n1816), .IN3(n353), .Q(n1815));
   XNOR3X1 U490 (.IN1(n838), .IN2(n1349), .IN3(n1350), .Q(n353));
   XNOR3X1 U491 (.IN1(n1346), .IN2(n1347), .IN3(n354), .Q(n1345));
   XNOR3X1 U492 (.IN1(n839), .IN2(n1349), .IN3(n1350), .Q(n354));
   XNOR3X1 U493 (.IN1(n508), .IN2(n618), .IN3(n355), .Q(n617));
   XNOR2X1 U494 (.IN1(n542), .IN2(n620), .Q(n355));
   INVX0 U495 (.INP(round_key[127]), .ZN(n1231));
   XNOR3X1 U496 (.IN1(n356), .IN2(n357), .IN3(n358), .Q(n1909));
   XNOR3X1 U497 (.IN1(n1531), .IN2(n1077), .IN3(n1913), .Q(n356));
   XNOR2X1 U498 (.IN1(n905), .IN2(n990), .Q(n357));
   XNOR3X1 U499 (.IN1(n1080), .IN2(n1078), .IN3(n1903), .Q(n358));
   INVX0 U500 (.INP(round_key[114]), .ZN(n1372));
   INVX0 U501 (.INP(round_key[19]), .ZN(n2193));
   XNOR2X1 U502 (.IN1(n930), .IN2(n999), .Q(n902));
   INVX0 U503 (.INP(round_key[83]), .ZN(n1719));
   XNOR3X1 U504 (.IN1(n667), .IN2(n740), .IN3(n359), .Q(n1702));
   XNOR2X1 U505 (.IN1(n742), .IN2(n634), .Q(n359));
   INVX0 U506 (.INP(n884), .ZN(n1809));
   XNOR2X1 U507 (.IN1(n984), .IN2(n360), .Q(n983));
   XNOR3X1 U508 (.IN1(n930), .IN2(n1614), .IN3(n986), .Q(n360));
   INVX0 U509 (.INP(n633), .ZN(n2207));
   INVX0 U510 (.INP(n1854), .ZN(n1634));
   INVX0 U511 (.INP(round_key[92]), .ZN(n1642));
   INVX0 U512 (.INP(n1184), .ZN(n2219));
   XNOR2X1 U513 (.IN1(n361), .IN2(n1624), .Q(n1622));
   XNOR3X1 U514 (.IN1(n639), .IN2(n740), .IN3(n1626), .Q(n361));
   XNOR2X1 U515 (.IN1(n362), .IN2(n632), .Q(n630));
   XNOR3X1 U516 (.IN1(n2183), .IN2(n636), .IN3(n637), .Q(n362));
   INVX0 U517 (.INP(n989), .ZN(n1892));
   XNOR2X1 U518 (.IN1(n1459), .IN2(n363), .Q(n1458));
   XNOR3X1 U519 (.IN1(n883), .IN2(n884), .IN3(n1461), .Q(n363));
   XNOR2X1 U520 (.IN1(n364), .IN2(n882), .Q(n880));
   XNOR3X1 U521 (.IN1(n1634), .IN2(n888), .IN3(n889), .Q(n364));
   XNOR3X1 U522 (.IN1(n365), .IN2(n366), .IN3(n367), .Q(n1389));
   XNOR2X1 U523 (.IN1(n778), .IN2(n776), .Q(n365));
   XNOR3X1 U524 (.IN1(n791), .IN2(n2169), .IN3(n772), .Q(n366));
   XNOR3X1 U525 (.IN1(n775), .IN2(n1393), .IN3(n774), .Q(n367));
   INVX0 U526 (.INP(n542), .ZN(n1348));
   XOR3X1 U527 (.IN1(n368), .IN2(n1529), .IN3(n369), .Q(n1527));
   XNOR2X1 U528 (.IN1(n1531), .IN2(n1075), .Q(n368));
   XNOR3X1 U529 (.IN1(n1080), .IN2(n1064), .IN3(n1863), .Q(n369));
   XNOR3X1 U530 (.IN1(n1179), .IN2(n370), .IN3(n1181), .Q(n1178));
   XNOR2X1 U531 (.IN1(n638), .IN2(n1184), .Q(n370));
   XNOR3X1 U532 (.IN1(n1841), .IN2(n371), .IN3(n1843), .Q(n1840));
   XNOR2X1 U533 (.IN1(n890), .IN2(n989), .Q(n371));
   XNOR3X1 U534 (.IN1(n1986), .IN2(n1987), .IN3(n372), .Q(n1985));
   XNOR3X1 U535 (.IN1(n990), .IN2(n1064), .IN3(n1863), .Q(n372));
   INVX0 U536 (.INP(n1714), .ZN(n2183));
   INVX0 U537 (.INP(round_key[28]), .ZN(n2184));
   XNOR2X1 U538 (.IN1(n373), .IN2(n585), .Q(n583));
   XOR3X1 U539 (.IN1(n589), .IN2(n590), .IN3(n591), .Q(n373));
   XNOR3X1 U540 (.IN1(n374), .IN2(n375), .IN3(n376), .Q(n1369));
   XNOR2X1 U541 (.IN1(n1373), .IN2(n870), .Q(n374));
   XNOR3X1 U542 (.IN1(n760), .IN2(n873), .IN3(n1314), .Q(n375));
   XOR3X1 U543 (.IN1(n750), .IN2(n861), .IN3(n854), .Q(n376));
   INVX0 U544 (.INP(round_key[113]), .ZN(n1377));
   INVX0 U545 (.INP(n578), .ZN(n1568));
   XNOR3X1 U546 (.IN1(n867), .IN2(n377), .IN3(n869), .Q(n866));
   XNOR2X1 U547 (.IN1(n750), .IN2(n767), .Q(n377));
   XNOR2X1 U548 (.IN1(n378), .IN2(n1383), .Q(n1381));
   XNOR3X1 U549 (.IN1(n761), .IN2(n809), .IN3(n1385), .Q(n378));
   XNOR3X1 U550 (.IN1(n1832), .IN2(n1833), .IN3(n379), .Q(n1831));
   XOR3X1 U551 (.IN1(n872), .IN2(n861), .IN3(n854), .Q(n379));
   INVX0 U552 (.INP(round_key[60]), .ZN(n1943));
   XNOR3X1 U553 (.IN1(n380), .IN2(n381), .IN3(n382), .Q(n1690));
   XNOR2X1 U554 (.IN1(n744), .IN2(n1279), .Q(n380));
   XNOR3X1 U555 (.IN1(n2181), .IN2(n743), .IN3(n1694), .Q(n381));
   XOR3X1 U556 (.IN1(n638), .IN2(n738), .IN3(n739), .Q(n382));
   XNOR3X1 U557 (.IN1(n734), .IN2(n735), .IN3(n383), .Q(n733));
   XOR3X1 U558 (.IN1(n737), .IN2(n738), .IN3(n739), .Q(n383));
   XNOR3X1 U559 (.IN1(n384), .IN2(n1927), .IN3(n1928), .Q(n1925));
   XNOR2X1 U560 (.IN1(n1399), .IN2(n557), .Q(n384));
   INVX0 U561 (.INP(round_key[51]), .ZN(n2150));
   XNOR3X1 U562 (.IN1(n1144), .IN2(n1145), .IN3(n385), .Q(n1143));
   XNOR3X1 U563 (.IN1(n592), .IN2(n1147), .IN3(n1148), .Q(n385));
   XNOR3X1 U564 (.IN1(n1144), .IN2(n1961), .IN3(n386), .Q(n1960));
   XNOR3X1 U565 (.IN1(n609), .IN2(n1147), .IN3(n1148), .Q(n386));
   INVX0 U566 (.INP(round_key[115]), .ZN(n1371));
   XNOR3X1 U567 (.IN1(n387), .IN2(n388), .IN3(n389), .Q(n1612));
   XNOR3X1 U568 (.IN1(n1173), .IN2(n621), .IN3(n1617), .Q(n387));
   XNOR2X1 U569 (.IN1(n516), .IN2(n547), .Q(n388));
   XNOR3X1 U570 (.IN1(n624), .IN2(n622), .IN3(n1416), .Q(n389));
   XNOR3X1 U571 (.IN1(n390), .IN2(n1170), .IN3(n1171), .Q(n1168));
   XNOR2X1 U572 (.IN1(n1173), .IN2(n620), .Q(n390));
   XNOR3X1 U573 (.IN1(n391), .IN2(n1978), .IN3(n1979), .Q(n1976));
   XNOR2X1 U574 (.IN1(n620), .IN2(n621), .Q(n391));
   XNOR3X1 U592 (.IN1(n392), .IN2(n393), .IN3(n394), .Q(n1273));
   XNOR3X1 U594 (.IN1(n743), .IN2(n1279), .IN3(n1280), .Q(n392));
   XNOR2X1 U596 (.IN1(n638), .IN2(n671), .Q(n393));
   XNOR3X1 U598 (.IN1(n737), .IN2(n1277), .IN3(n1278), .Q(n394));
   INVX0 U600 (.INP(n809), .ZN(n2149));
   XNOR3X1 U602 (.IN1(n395), .IN2(n396), .IN3(n397), .Q(n1769));
   XNOR2X1 U604 (.IN1(n775), .IN2(n875), .Q(n395));
   XNOR3X1 U606 (.IN1(n808), .IN2(n760), .IN3(n1773), .Q(n396));
   XNOR3X1 U608 (.IN1(n750), .IN2(n1289), .IN3(n1290), .Q(n397));
   XNOR3X1 U610 (.IN1(n398), .IN2(n399), .IN3(n400), .Q(n1285));
   XNOR2X1 U612 (.IN1(n875), .IN2(n1912), .Q(n398));
   XNOR3X1 U614 (.IN1(n808), .IN2(n760), .IN3(n1291), .Q(n399));
   XNOR3X1 U641 (.IN1(n751), .IN2(n1289), .IN3(n1290), .Q(n400));
   INVX0 U644 (.INP(n755), .ZN(n2173));
   INVX0 U650 (.INP(n517), .ZN(n1549));
   XNOR2X1 U652 (.IN1(n401), .IN2(n507), .Q(n504));
   XNOR3X1 U658 (.IN1(n513), .IN2(n514), .IN3(n515), .Q(n401));
   XNOR3X1 U659 (.IN1(n402), .IN2(n403), .IN3(n404), .Q(n1536));
   XNOR3X1 U667 (.IN1(n1093), .IN2(n618), .IN3(n1541), .Q(n402));
   XNOR2X1 U670 (.IN1(n516), .IN2(n517), .Q(n403));
   XNOR3X1 U676 (.IN1(n513), .IN2(n514), .IN3(n1540), .Q(n404));
   INVX0 U679 (.INP(n601), .ZN(n1497));
   INVX0 U685 (.INP(n514), .ZN(n1370));
   XNOR3X1 U687 (.IN1(n405), .IN2(n406), .IN3(n407), .Q(n1086));
   XNOR2X1 U693 (.IN1(n1093), .IN2(n618), .Q(n405));
   XNOR3X1 U696 (.IN1(n509), .IN2(n540), .IN3(n1092), .Q(n406));
   XNOR3X1 U703 (.IN1(n516), .IN2(n1090), .IN3(n1091), .Q(n407));
   XNOR3X1 U704 (.IN1(n1597), .IN2(n408), .IN3(n1920), .Q(n1918));
   XNOR3X1 U711 (.IN1(n508), .IN2(n540), .IN3(n1092), .Q(n408));
   INVX0 U713 (.INP(round_key[124]), .ZN(n1263));
   INVX0 U718 (.INP(round_key[52]), .ZN(n2148));
   INVX0 U721 (.INP(round_key[76]), .ZN(n1801));
   INVX0 U726 (.INP(round_key[44]), .ZN(n2161));
   INVX0 U727 (.INP(round_key[12]), .ZN(n2206));
   INVX0 U734 (.INP(round_key[84]), .ZN(n1709));
   INVX0 U736 (.INP(round_key[20]), .ZN(n2192));
   INVX0 U743 (.INP(round_key[36]), .ZN(n2172));
   INVX0 U744 (.INP(round_key[100]), .ZN(n1548));
   INVX0 U748 (.INP(round_key[105]), .ZN(n1486));
   INVX0 U749 (.INP(round_key[99]), .ZN(n1556));
   INVX0 U757 (.INP(round_key[68]), .ZN(n1883));
   INVX0 U758 (.INP(round_key[4]), .ZN(n2218));
   INVX0 U762 (.INP(round_key[3]), .ZN(n2220));
   INVX0 U763 (.INP(round_key[35]), .ZN(n2174));
   INVX0 U771 (.INP(round_key[87]), .ZN(n1691));
   INVX0 U774 (.INP(round_key[79]), .ZN(n1752));
   INVX0 U778 (.INP(round_key[15]), .ZN(n2197));
   INVX0 U779 (.INP(round_key[77]), .ZN(n1779));
   INVX0 U787 (.INP(round_key[46]), .ZN(n2157));
   INVX0 U788 (.INP(round_key[45]), .ZN(n2160));
   INVX0 U790 (.INP(round_key[55]), .ZN(n1988));
   INVX0 U794 (.INP(round_key[78]), .ZN(n1770));
   INVX0 U796 (.INP(round_key[53]), .ZN(n2146));
   INVX0 U802 (.INP(round_key[14]), .ZN(n2201));
   INVX0 U804 (.INP(round_key[85]), .ZN(n1696));
   INVX0 U810 (.INP(round_key[54]), .ZN(n2144));
   INVX0 U811 (.INP(round_key[13]), .ZN(n2204));
   INVX0 U812 (.INP(round_key[86]), .ZN(n1692));
   INVX0 U813 (.INP(round_key[47]), .ZN(n2154));
   INVX0 U818 (.INP(round_key[103]), .ZN(n1528));
   INVX0 U821 (.INP(round_key[7]), .ZN(n2212));
   INVX0 U826 (.INP(round_key[39]), .ZN(n2166));
   INVX0 U828 (.INP(round_key[101]), .ZN(n1538));
   INVX0 U834 (.INP(round_key[102]), .ZN(n1530));
   INVX0 U837 (.INP(round_key[71]), .ZN(n1852));
   INVX0 U842 (.INP(round_key[37]), .ZN(n2170));
   INVX0 U845 (.INP(round_key[6]), .ZN(n2214));
   INVX0 U850 (.INP(round_key[70]), .ZN(n1862));
   INVX0 U851 (.INP(round_key[5]), .ZN(n2216));
   INVX0 U856 (.INP(round_key[69]), .ZN(n1871));
   INVX0 U857 (.INP(round_key[38]), .ZN(n2168));
   INVX0 U863 (.INP(round_key[56]), .ZN(n1977));
   INVX0 U864 (.INP(round_key[63]), .ZN(n1911));
   INVX0 U877 (.INP(round_key[95]), .ZN(n1606));
   INVX0 U878 (.INP(round_key[58]), .ZN(n1962));
   INVX0 U884 (.INP(round_key[90]), .ZN(n1661));
   INVX0 U885 (.INP(round_key[91]), .ZN(n1651));
   INVX0 U893 (.INP(round_key[89]), .ZN(n1674));
   INVX0 U896 (.INP(round_key[25]), .ZN(n2187));
   INVX0 U902 (.INP(round_key[59]), .ZN(n1953));
   INVX0 U905 (.INP(round_key[57]), .ZN(n1970));
   INVX0 U911 (.INP(round_key[88]), .ZN(n1682));
   INVX0 U912 (.INP(round_key[31]), .ZN(n2179));
   INVX0 U920 (.INP(round_key[27]), .ZN(n2185));
   INVX0 U923 (.INP(round_key[26]), .ZN(n2186));
   INVX0 U929 (.INP(round_key[24]), .ZN(n2188));
   INVX0 U932 (.INP(round_key[116]), .ZN(n1360));
   INVX0 U938 (.INP(round_key[108]), .ZN(n1460));
   INVX0 U941 (.INP(round_key[111]), .ZN(n1390));
   INVX0 U948 (.INP(round_key[119]), .ZN(n1287));
   INVX0 U949 (.INP(round_key[117]), .ZN(n1324));
   INVX0 U956 (.INP(round_key[110]), .ZN(n1407));
   INVX0 U957 (.INP(round_key[118]), .ZN(n1297));
   INVX0 U958 (.INP(round_key[109]), .ZN(n1450));
   OA21X1 U959 (.IN1(round_key[20]), .IN2(n440), .IN3(n457), .Q(n1794));
   OA21X1 U963 (.IN1(round_key[105]), .IN2(n519), .IN3(n625), .Q(n847));
   OA21X1 U965 (.IN1(round_key[36]), .IN2(n444), .IN3(n1453), .Q(n1647));
   OA21X1 U967 (.IN1(round_key[12]), .IN2(n897), .IN3(n457), .Q(n1867));
   OA21X1 U971 (.IN1(round_key[52]), .IN2(n440), .IN3(n462), .Q(n1483));
   OA21X1 U972 (.IN1(round_key[44]), .IN2(n868), .IN3(n462), .Q(n1565));
   OA21X1 U979 (.IN1(round_key[76]), .IN2(n881), .IN3(n538), .Q(n1213));
   OA21X1 U980 (.IN1(round_key[84]), .IN2(n443), .IN3(n538), .Q(n1117));
   OA21X1 U984 (.IN1(round_key[4]), .IN2(n868), .IN3(n458), .Q(n1939));
   OA21X1 U985 (.IN1(round_key[99]), .IN2(n446), .IN3(n625), .Q(n934));
   OA21X1 U991 (.IN1(round_key[100]), .IN2(n445), .IN3(n625), .Q(n921));
   OA21X1 U992 (.IN1(round_key[35]), .IN2(n448), .IN3(n1453), .Q(n1657));
   OA21X1 U1005 (.IN1(round_key[3]), .IN2(n445), .IN3(n458), .Q(n1949));
   OA21X1 U1009 (.IN1(round_key[68]), .IN2(n445), .IN3(n553), .Q(n1319));
   OA21X1 U1013 (.IN1(round_key[45]), .IN2(n850), .IN3(n462), .Q(n1553));
   OA21X1 U1015 (.IN1(round_key[15]), .IN2(n441), .IN3(n457), .Q(n1838));
   OA21X1 U1021 (.IN1(round_key[71]), .IN2(n850), .IN3(n553), .Q(n1283));
   OA21X1 U1022 (.IN1(round_key[87]), .IN2(n850), .IN3(n538), .Q(n1084));
   OA21X1 U1023 (.IN1(round_key[79]), .IN2(n438), .IN3(n538), .Q(n1176));
   OA21X1 U1029 (.IN1(round_key[53]), .IN2(n897), .IN3(n462), .Q(n1474));
   OA21X1 U1030 (.IN1(round_key[55]), .IN2(n445), .IN3(n462), .Q(n1456));
   OA21X1 U1032 (.IN1(round_key[54]), .IN2(n445), .IN3(n462), .Q(n1465));
   OA21X1 U1033 (.IN1(round_key[47]), .IN2(n440), .IN3(n462), .Q(n1534));
   OA21X1 U1037 (.IN1(round_key[14]), .IN2(n850), .IN3(n457), .Q(n1847));
   OA21X1 U1038 (.IN1(round_key[13]), .IN2(n439), .IN3(n457), .Q(n1858));
   OA21X1 U1039 (.IN1(round_key[101]), .IN2(n897), .IN3(n625), .Q(n909));
   OA21X1 U1040 (.IN1(round_key[86]), .IN2(n436), .IN3(n538), .Q(n1096));
   OA21X1 U1045 (.IN1(round_key[77]), .IN2(n448), .IN3(n538), .Q(n1200));
   OA21X1 U1047 (.IN1(round_key[46]), .IN2(n448), .IN3(n462), .Q(n1544));
   OA21X1 U1053 (.IN1(round_key[78]), .IN2(n438), .IN3(n538), .Q(n1188));
   OA21X1 U1055 (.IN1(round_key[85]), .IN2(n440), .IN3(n538), .Q(n1107));
   OA21X1 U1056 (.IN1(round_key[103]), .IN2(n881), .IN3(n625), .Q(n878));
   OA21X1 U1061 (.IN1(round_key[39]), .IN2(n442), .IN3(n1453), .Q(n1620));
   OA21X1 U1062 (.IN1(round_key[6]), .IN2(n447), .IN3(n458), .Q(n1923));
   OA21X1 U1063 (.IN1(round_key[7]), .IN2(n448), .IN3(n458), .Q(n1916));
   OA21X1 U1064 (.IN1(round_key[69]), .IN2(n444), .IN3(n553), .Q(n1306));
   OA21X1 U1069 (.IN1(round_key[5]), .IN2(n446), .IN3(n458), .Q(n1931));
   OA21X1 U1070 (.IN1(round_key[38]), .IN2(n443), .IN3(n1453), .Q(n1629));
   OA21X1 U1071 (.IN1(round_key[37]), .IN2(n443), .IN3(n1453), .Q(n1638));
   OA21X1 U1072 (.IN1(round_key[70]), .IN2(n868), .IN3(n553), .Q(n1294));
   OA21X1 U1077 (.IN1(round_key[102]), .IN2(n444), .IN3(n625), .Q(n894));
   OA21X1 U1078 (.IN1(round_key[49]), .IN2(n436), .IN3(n462), .Q(n1516));
   OA21X1 U1079 (.IN1(round_key[19]), .IN2(n446), .IN3(n457), .Q(n1804));
   OA21X1 U1081 (.IN1(round_key[43]), .IN2(n439), .IN3(n462), .Q(n1576));
   OA21X1 U1085 (.IN1(round_key[65]), .IN2(n850), .IN3(n553), .Q(n1355));
   OA21X1 U1089 (.IN1(round_key[17]), .IN2(n897), .IN3(n457), .Q(n1821));
   OA21X1 U1093 (.IN1(round_key[81]), .IN2(n445), .IN3(n538), .Q(n1153));
   OA21X1 U1095 (.IN1(round_key[83]), .IN2(n444), .IN3(n538), .Q(n1128));
   OA21X1 U1100 (.IN1(round_key[51]), .IN2(n850), .IN3(n462), .Q(n1493));
   OA21X1 U1101 (.IN1(round_key[11]), .IN2(n868), .IN3(n457), .Q(n1879));
   OA21X1 U1114 (.IN1(round_key[75]), .IN2(n439), .IN3(n538), .Q(n1227));
   OA21X1 U1115 (.IN1(round_key[67]), .IN2(n445), .IN3(n553), .Q(n1330));
   OA21X1 U1121 (.IN1(round_key[1]), .IN2(n881), .IN3(n458), .Q(n1966));
   OA21X1 U1122 (.IN1(round_key[41]), .IN2(n519), .IN3(n1453), .Q(n1601));
   OA21X1 U1128 (.IN1(round_key[73]), .IN2(n881), .IN3(n553), .Q(n1258));
   OA21X1 U1129 (.IN1(round_key[97]), .IN2(n448), .IN3(n625), .Q(n966));
   OA21X1 U1130 (.IN1(round_key[9]), .IN2(n436), .IN3(n458), .Q(n1897));
   OA21X1 U1132 (.IN1(round_key[33]), .IN2(n442), .IN3(n1453), .Q(n1679));
   OA21X1 U1134 (.IN1(round_key[23]), .IN2(n441), .IN3(n457), .Q(n1767));
   OA21X1 U1137 (.IN1(round_key[80]), .IN2(n439), .IN3(n538), .Q(n1166));
   OA21X1 U1140 (.IN1(round_key[48]), .IN2(n444), .IN3(n462), .Q(n1525));
   OA21X1 U1147 (.IN1(round_key[22]), .IN2(n442), .IN3(n457), .Q(n1776));
   OA21X1 U1148 (.IN1(round_key[66]), .IN2(n446), .IN3(n553), .Q(n1343));
   OA21X1 U1149 (.IN1(round_key[8]), .IN2(n881), .IN3(n458), .Q(n1907));
   OA21X1 U1151 (.IN1(round_key[40]), .IN2(n441), .IN3(n1453), .Q(n1610));
   OA21X1 U1152 (.IN1(round_key[72]), .IN2(n441), .IN3(n553), .Q(n1271));
   OA21X1 U1158 (.IN1(round_key[64]), .IN2(n447), .IN3(n553), .Q(n1367));
   OA21X1 U1159 (.IN1(round_key[18]), .IN2(n438), .IN3(n457), .Q(n1813));
   OA21X1 U1169 (.IN1(round_key[32]), .IN2(n443), .IN3(n1453), .Q(n1688));
   OA21X1 U1170 (.IN1(round_key[21]), .IN2(n439), .IN3(n457), .Q(n1785));
   OA21X1 U1180 (.IN1(round_key[16]), .IN2(n447), .IN3(n457), .Q(n1829));
   OA21X1 U1183 (.IN1(round_key[50]), .IN2(n439), .IN3(n462), .Q(n1506));
   OA21X1 U1202 (.IN1(round_key[82]), .IN2(n438), .IN3(n538), .Q(n1141));
   OA21X1 U1203 (.IN1(round_key[104]), .IN2(n439), .IN3(n625), .Q(n864));
   OA21X1 U1214 (.IN1(round_key[2]), .IN2(n897), .IN3(n458), .Q(n1958));
   OA21X1 U1215 (.IN1(round_key[74]), .IN2(n442), .IN3(n553), .Q(n1244));
   OA21X1 U1222 (.IN1(round_key[42]), .IN2(n440), .IN3(n1453), .Q(n1590));
   OA21X1 U1223 (.IN1(round_key[10]), .IN2(n447), .IN3(n458), .Q(n1888));
   OA21X1 U1233 (.IN1(round_key[96]), .IN2(n438), .IN3(n625), .Q(n1983));
   OA21X1 U1234 (.IN1(round_key[34]), .IN2(n444), .IN3(n1453), .Q(n1670));
   OA21X1 U1238 (.IN1(round_key[0]), .IN2(n441), .IN3(n458), .Q(n1974));
   OA21X1 U1242 (.IN1(round_key[106]), .IN2(n446), .IN3(n625), .Q(n829));
   OA21X1 U1246 (.IN1(round_key[98]), .IN2(n447), .IN3(n625), .Q(n950));
   INVX0 U1247 (.INP(round_key[120]), .ZN(n1286));
   INVX0 U1251 (.INP(round_key[121]), .ZN(n1276));
   INVX0 U1253 (.INP(round_key[123]), .ZN(n1274));
   INVX0 U1254 (.INP(round_key[122]), .ZN(n1275));
   AND2X1 U1255 (.IN1(n1375), .IN2(n497), .Q(n409));
   NAND2X1 U1261 (.IN1(n1994), .IN2(n2001), .QN(n2139));
   INVX0 U1262 (.INP(n1994), .ZN(n2230));
   NAND2X1 U1281 (.IN1(n2229), .IN2(n1980), .QN(n2001));
   INVX0 U1282 (.INP(n1993), .ZN(n2229));
   NAND2X1 U1291 (.IN1(n833), .IN2(n315), .QN(n782));
   NAND2X1 U1292 (.IN1(n435), .IN2(n272), .QN(n1201));
   NAND2X1 U1295 (.IN1(n834), .IN2(n300), .QN(n661));
   NAND2X1 U1299 (.IN1(n834), .IN2(n239), .QN(n1639));
   NAND2X1 U1300 (.IN1(n914), .IN2(n302), .QN(n676));
   NAND2X1 U1304 (.IN1(n914), .IN2(n241), .QN(n1648));
   NAND2X1 U1305 (.IN1(n816), .IN2(n215), .QN(n1484));
   NAND2X1 U1310 (.IN1(n833), .IN2(n330), .QN(n922));
   NAND2X1 U1311 (.IN1(n833), .IN2(n313), .QN(n765));
   NAND2X1 U1312 (.IN1(n832), .IN2(n298), .QN(n644));
   NAND2X1 U1314 (.IN1(n834), .IN2(n317), .QN(n797));
   NAND2X1 U1319 (.IN1(n816), .IN2(n274), .QN(n1214));
   NAND2X1 U1320 (.IN1(n914), .IN2(n318), .QN(n813));
   NAND2X0 U1329 (.IN1(n437), .IN2(n303), .QN(n688));
   NAND2X1 U1330 (.IN1(n914), .IN2(n225), .QN(n1545));
   NAND2X1 U1339 (.IN1(n435), .IN2(n229), .QN(n1566));
   NAND2X1 U1340 (.IN1(n434), .IN2(n227), .QN(n1554));
   NAND2X1 U1350 (.IN1(n832), .IN2(n243), .QN(n1658));
   NAND2X1 U1351 (.IN1(n832), .IN2(n275), .QN(n1228));
   NAND2X0 U1354 (.IN1(n434), .IN2(n185), .QN(n1880));
   NAND2X1 U1360 (.IN1(n434), .IN2(n218), .QN(n1517));
   NAND2X1 U1364 (.IN1(n816), .IN2(n334), .QN(n967));
   NAND2X0 U1369 (.IN1(n437), .IN2(n216), .QN(n1494));
   NAND2X1 U1370 (.IN1(n914), .IN2(n332), .QN(n935));
   NAND2X1 U1371 (.IN1(n914), .IN2(n169), .QN(n1795));
   NAND2X1 U1372 (.IN1(n435), .IN2(n288), .QN(n1320));
   NAND2X0 U1377 (.IN1(n833), .IN2(n213), .QN(n1475));
   NAND2X1 U1381 (.IN1(n786), .IN2(n328), .QN(n910));
   NAND2X1 U1387 (.IN1(n786), .IN2(n197), .QN(n1940));
   NAND2X1 U1388 (.IN1(n435), .IN2(n187), .QN(n1898));
   NAND2X0 U1392 (.IN1(n435), .IN2(n186), .QN(n1889));
   NAND2X1 U1393 (.IN1(n434), .IN2(n167), .QN(n1786));
   NAND2X1 U1397 (.IN1(n832), .IN2(n286), .QN(n1307));
   NAND2X1 U1398 (.IN1(n800), .IN2(n170), .QN(n1805));
   NAND2X1 U1406 (.IN1(n833), .IN2(n230), .QN(n1577));
   NAND2X0 U1407 (.IN1(n435), .IN2(n260), .QN(n1118));
   NAND2X1 U1408 (.IN1(n786), .IN2(n184), .QN(n1868));
   NAND2X0 U1409 (.IN1(n816), .IN2(n211), .QN(n1466));
   NAND2X1 U1416 (.IN1(n834), .IN2(n326), .QN(n895));
   NAND2X0 U1417 (.IN1(n832), .IN2(n232), .QN(n1602));
   NAND2X1 U1426 (.IN1(n816), .IN2(n291), .QN(n1356));
   NAND2X0 U1427 (.IN1(n435), .IN2(n172), .QN(n1822));
   NAND2X0 U1436 (.IN1(n800), .IN2(n277), .QN(n1259));
   NAND2X0 U1440 (.IN1(n437), .IN2(n258), .QN(n1108));
   NAND2X0 U1446 (.IN1(n914), .IN2(n195), .QN(n1932));
   NAND2X0 U1447 (.IN1(n437), .IN2(n321), .QN(n848));
   NAND2X1 U1448 (.IN1(n786), .IN2(n305), .QN(n718));
   NAND2X0 U1450 (.IN1(n914), .IN2(n245), .QN(n1680));
   NAND2X0 U1452 (.IN1(n816), .IN2(n319), .QN(n830));
   NAND2X1 U1456 (.IN1(n434), .IN2(n237), .QN(n1630));
   NAND2X0 U1457 (.IN1(n435), .IN2(n166), .QN(n1777));
   NAND2X0 U1466 (.IN1(n832), .IN2(n284), .QN(n1295));
   NAND2X0 U1469 (.IN1(n786), .IN2(n289), .QN(n1331));
   NAND2X1 U1478 (.IN1(n800), .IN2(n307), .QN(n748));
   NAND2X0 U1482 (.IN1(n816), .IN2(n231), .QN(n1591));
   NAND2X0 U1494 (.IN1(n833), .IN2(n182), .QN(n1859));
   NAND2X0 U1502 (.IN1(n832), .IN2(n256), .QN(n1097));
   NAND2X0 U1521 (.IN1(n834), .IN2(n180), .QN(n1848));
   NAND2X0 U1522 (.IN1(n834), .IN2(n270), .QN(n1189));
   NAND2X0 U1537 (.IN1(n434), .IN2(n261), .QN(n1129));
   NAND2X0 U1544 (.IN1(n437), .IN2(n199), .QN(n1950));
   NAND2X1 U1550 (.IN1(n800), .IN2(n304), .QN(n702));
   NAND2X0 U1563 (.IN1(n434), .IN2(n244), .QN(n1671));
   NAND2X0 U1571 (.IN1(n833), .IN2(n201), .QN(n1967));
   NAND2X0 U1582 (.IN1(n914), .IN2(n263), .QN(n1154));
   NAND2X0 U1587 (.IN1(n434), .IN2(n276), .QN(n1245));
   NAND2X0 U1591 (.IN1(n914), .IN2(n171), .QN(n1814));
   NAND2X1 U1593 (.IN1(n800), .IN2(n290), .QN(n1344));
   NAND2X0 U1594 (.IN1(n434), .IN2(n188), .QN(n1908));
   NAND2X0 U1609 (.IN1(n435), .IN2(n217), .QN(n1507));
   NAND2X0 U1610 (.IN1(n833), .IN2(n333), .QN(n951));
   NAND2X0 U1613 (.IN1(n834), .IN2(n234), .QN(n1621));
   NAND2X0 U1615 (.IN1(n800), .IN2(n296), .QN(n629));
   NAND2X0 U1619 (.IN1(n435), .IN2(n209), .QN(n1457));
   NAND2X0 U1626 (.IN1(n800), .IN2(n323), .QN(n879));
   NAND2X0 U1630 (.IN1(n786), .IN2(n219), .QN(n1526));
   NAND2X0 U1638 (.IN1(n786), .IN2(n265), .QN(n1177));
   NAND2X0 U1655 (.IN1(n816), .IN2(n177), .QN(n1839));
   NAND2X0 U1656 (.IN1(n786), .IN2(n335), .QN(n1984));
   NAND2X0 U1679 (.IN1(n914), .IN2(n292), .QN(n1368));
   NAND2X0 U1680 (.IN1(n833), .IN2(n322), .QN(n865));
   NAND2X0 U1687 (.IN1(n914), .IN2(n173), .QN(n1830));
   NAND2X0 U1693 (.IN1(n834), .IN2(n306), .QN(n732));
   NAND2X0 U1694 (.IN1(n434), .IN2(n246), .QN(n1689));
   NAND2X0 U1719 (.IN1(n800), .IN2(n193), .QN(n1924));
   NAND2X0 U1720 (.IN1(n834), .IN2(n262), .QN(n1142));
   NAND2X0 U1734 (.IN1(n816), .IN2(n200), .QN(n1959));
   NAND2X0 U1735 (.IN1(n832), .IN2(n233), .QN(n1611));
   NAND2X0 U1755 (.IN1(n437), .IN2(n264), .QN(n1167));
   NAND2X0 U1759 (.IN1(n786), .IN2(n202), .QN(n1975));
   NAND2X0 U1765 (.IN1(n437), .IN2(n278), .QN(n1272));
   NAND2X0 U1766 (.IN1(n786), .IN2(n164), .QN(n1768));
   NAND2X0 U1776 (.IN1(n832), .IN2(n280), .QN(n1284));
   NAND2X0 U1777 (.IN1(n435), .IN2(n222), .QN(n1535));
   NAND2X0 U1782 (.IN1(n437), .IN2(n253), .QN(n1085));
   NAND2X0 U1783 (.IN1(n914), .IN2(n190), .QN(n1917));
   AO22X1 U1791 (.IN1(new_block[117]), .IN2(n454), .IN3(new_block[85]), .IN4(n449), .Q(
          n482));
   NOR4X0 U1792 (.IN1(round[0]), .IN2(round[1]), .IN3(round[2]), .IN4(round[3]), .QN(n1992)
          );
   NAND2X0 U1802 (.IN1(dec_ctrl_reg[1]), .IN2(n159), .QN(n1993));
   NAND3X0 U1805 (.IN1(n159), .IN2(n158), .IN3(next), .QN(n1994));
   NOR2X0 U1816 (.IN1(n205), .IN2(sword_ctr_reg[1]), .QN(n1376));
   NOR2X0 U1822 (.IN1(n204), .IN2(n205), .QN(n1980));
   NOR2X0 U1825 (.IN1(n204), .IN2(sword_ctr_reg[0]), .QN(n1695));
   NOR2X0 U1839 (.IN1(round[2]), .IN2(round[1]), .QN(n1998));
   AO22X1 U1845 (.IN1(new_block[125]), .IN2(n454), .IN3(new_block[93]), .IN4(n450), .Q(
          n474));
   AO22X1 U1857 (.IN1(new_block[120]), .IN2(n454), .IN3(new_block[88]), .IN4(n450), .Q(
          n479));
   AO22X1 U1858 (.IN1(new_block[121]), .IN2(n454), .IN3(new_block[89]), .IN4(n450), .Q(
          n478));
   AO22X1 U1863 (.IN1(new_block[124]), .IN2(n454), .IN3(new_block[92]), .IN4(n449), .Q(
          n475));
   AO22X1 U1866 (.IN1(new_block[116]), .IN2(n454), .IN3(new_block[84]), .IN4(n450), .Q(
          n483));
   AO22X1 U1874 (.IN1(new_block[123]), .IN2(n454), .IN3(new_block[91]), .IN4(n449), .Q(
          n476));
   AO22X1 U1875 (.IN1(new_block[122]), .IN2(n454), .IN3(new_block[90]), .IN4(n450), .Q(
          n477));
   AO22X1 U1881 (.IN1(new_block[98]), .IN2(n454), .IN3(new_block[66]), .IN4(n450), .Q(n473)
          );
   AO22X1 U1882 (.IN1(new_block[118]), .IN2(n454), .IN3(new_block[86]), .IN4(n450), .Q(
          n481));
   AO22X1 U1888 (.IN1(new_block[126]), .IN2(n454), .IN3(new_block[94]), .IN4(n449), .Q(
          n472));
   AO22X1 U1892 (.IN1(new_block[119]), .IN2(n454), .IN3(new_block[87]), .IN4(n450), .Q(
          n480));
   NOR2X0 U1897 (.IN1(n2001), .IN2(round[0]), .QN(n1999));
   NBUFFX2 U2074 (.INP(n897), .Z(n448));
   NBUFFX2 U2075 (.INP(n897), .Z(n447));
   NBUFFX2 U2076 (.INP(n897), .Z(n446));
   NBUFFX2 U2077 (.INP(n448), .Z(n438));
   NBUFFX2 U2078 (.INP(n448), .Z(n439));
   NBUFFX2 U2079 (.INP(n446), .Z(n445));
   NBUFFX2 U2080 (.INP(n446), .Z(n444));
   NBUFFX2 U2081 (.INP(n447), .Z(n440));
   NBUFFX2 U2082 (.INP(n447), .Z(n441));
   NBUFFX2 U2083 (.INP(n447), .Z(n442));
   NBUFFX2 U2084 (.INP(n446), .Z(n443));
   INVX0 U2085 (.INP(n437), .ZN(n436));
   INVX0 U2086 (.INP(n881), .ZN(n437));
   INVX0 U2087 (.INP(n850), .ZN(n434));
   INVX0 U2088 (.INP(n868), .ZN(n435));
   INVX0 U2089 (.INP(n499), .ZN(n451));
   INVX0 U2090 (.INP(n496), .ZN(n449));
   INVX0 U2091 (.INP(n496), .ZN(n450));
   INVX0 U2092 (.INP(n499), .ZN(n452));
   INVX0 U2093 (.INP(n463), .ZN(n462));
   INVX0 U2094 (.INP(n1453), .ZN(n463));
   OA21X1 U2095 (.IN1(n2228), .IN2(n1992), .IN3(n2003), .Q(n1990));
   INVX0 U2096 (.INP(n1995), .ZN(n2228));
   INVX0 U2097 (.INP(n1990), .ZN(n2227));
   NOR2X0 U2098 (.IN1(n2227), .IN2(n1991), .QN(n1374));
   INVX0 U2099 (.INP(n142), .ZN(n506));
   INVX0 U2100 (.INP(n142), .ZN(n500));
   INVX0 U2101 (.INP(n142), .ZN(n525));
   INVX0 U2102 (.INP(n753), .ZN(n736));
   INVX0 U2103 (.INP(n753), .ZN(n706));
   INVX0 U2104 (.INP(n753), .ZN(n727));
   INVX0 U2105 (.INP(n753), .ZN(n631));
   INVX0 U2106 (.INP(n753), .ZN(n646));
   INVX0 U2107 (.INP(n753), .ZN(n664));
   INVX0 U2108 (.INP(n753), .ZN(n679));
   INVX0 U2109 (.INP(n753), .ZN(n697));
   INVX0 U2110 (.INP(n4), .ZN(n584));
   INVX0 U2111 (.INP(n4), .ZN(n567));
   INVX0 U2112 (.INP(n4), .ZN(n599));
   NAND2X0 U2113 (.IN1(n1695), .IN2(n1374), .QN(n498));
   NAND2X0 U2114 (.IN1(n1980), .IN2(n1374), .QN(n499));
   OA21X1 U2115 (.IN1(round_key[113]), .IN2(n519), .IN3(n619), .Q(n717));
   OA21X1 U2116 (.IN1(round_key[117]), .IN2(n868), .IN3(n619), .Q(n660));
   OA21X1 U2117 (.IN1(round_key[108]), .IN2(n519), .IN3(n619), .Q(n796));
   OA21X1 U2118 (.IN1(round_key[111]), .IN2(n441), .IN3(n619), .Q(n747));
   OA21X1 U2119 (.IN1(round_key[115]), .IN2(n440), .IN3(n619), .Q(n687));
   OA21X1 U2120 (.IN1(round_key[114]), .IN2(n850), .IN3(n619), .Q(n701));
   OA21X1 U2121 (.IN1(round_key[112]), .IN2(n447), .IN3(n619), .Q(n731));
   OA21X1 U2122 (.IN1(round_key[107]), .IN2(n441), .IN3(n619), .Q(n812));
   OA21X1 U2123 (.IN1(round_key[119]), .IN2(n436), .IN3(n619), .Q(n628));
   OA21X1 U2124 (.IN1(round_key[118]), .IN2(n868), .IN3(n619), .Q(n643));
   OA21X1 U2125 (.IN1(round_key[116]), .IN2(n519), .IN3(n619), .Q(n675));
   OA21X1 U2126 (.IN1(round_key[110]), .IN2(n868), .IN3(n619), .Q(n764));
   OA21X1 U2127 (.IN1(round_key[109]), .IN2(n444), .IN3(n619), .Q(n781));
   INVX0 U2128 (.INP(n497), .ZN(n454));
   INVX0 U2129 (.INP(n497), .ZN(n453));
   INVX0 U2130 (.INP(n800), .ZN(n897));
   INVX0 U2131 (.INP(n914), .ZN(n850));
   INVX0 U2132 (.INP(n914), .ZN(n868));
   INVX0 U2133 (.INP(n519), .ZN(n914));
   INVX0 U2134 (.INP(n850), .ZN(n834));
   INVX0 U2135 (.INP(n850), .ZN(n832));
   INVX0 U2136 (.INP(n850), .ZN(n833));
   INVX0 U2137 (.INP(n868), .ZN(n786));
   INVX0 U2138 (.INP(n868), .ZN(n800));
   INVX0 U2139 (.INP(n868), .ZN(n816));
   INVX0 U2140 (.INP(n1), .ZN(n553));
   INVX0 U2141 (.INP(n409), .ZN(n625));
   INVX0 U2142 (.INP(n498), .ZN(n455));
   NAND2X0 U2143 (.IN1(dec_ctrl_reg[0]), .IN2(n158), .QN(n2003));
   NAND2X0 U2144 (.IN1(n1376), .IN2(n1374), .QN(n496));
   INVX0 U2145 (.INP(n144), .ZN(n457));
   INVX0 U2146 (.INP(n144), .ZN(n458));
   INVX0 U2147 (.INP(n3), .ZN(n461));
   NAND2X0 U2148 (.IN1(n1375), .IN2(n498), .QN(n1453));
   NOR2X0 U2149 (.IN1(n158), .IN2(n159), .QN(n1995));
   INVX0 U2150 (.INP(n3), .ZN(n459));
   INVX0 U2151 (.INP(n3), .ZN(n460));
   OA21X1 U2152 (.IN1(n2228), .IN2(n1992), .IN3(n1993), .Q(n1991));
   INVX0 U2153 (.INP(n409), .ZN(n619));
   INVX0 U2154 (.INP(n1), .ZN(n538));
   INVX0 U2155 (.INP(n914), .ZN(n881));
   NAND2X0 U2156 (.IN1(n1992), .IN2(n1995), .QN(n519));
   INVX0 U2157 (.INP(n785), .ZN(n753));
   INVX0 U2158 (.INP(n785), .ZN(n768));
   INVX0 U2159 (.INP(n520), .ZN(n785));
   NAND2X0 U2160 (.IN1(n1991), .IN2(n2227), .QN(n520));
   XOR2X2 U2161 (.IN1(n164), .IN2(n2189), .Q(n740));
   XOR2X2 U2162 (.IN1(n167), .IN2(n2191), .Q(n649));
   XOR2X2 U2163 (.IN1(n166), .IN2(n2190), .Q(n634));
endmodule

module aes_key_mem_test_1 (clk, reset_n, key, keylen, init, round, round_key, ready, sboxw
       , new_sboxw, test_si3, test_si2, test_si1, test_so3, test_so2, test_so1, test_se);
input clk, reset_n, keylen, init, test_si3, test_si2, test_si1, test_se;
input [255:0] key;
input [3:0] round;
input [31:0] new_sboxw;
output ready, test_so3, test_so2, test_so1;
output [127:0] round_key;
output [31:0] sboxw;
wire N28, N29, N30, N31, \key_mem[0][127] , \key_mem[0][126] , \key_mem[0][125] , 
       \key_mem[0][124] , \key_mem[0][123] , \key_mem[0][122] , \key_mem[0][121] , 
       \key_mem[0][120] , \key_mem[0][119] , \key_mem[0][118] , \key_mem[0][117] , 
       \key_mem[0][116] , \key_mem[0][115] , \key_mem[0][114] , \key_mem[0][113] , 
       \key_mem[0][112] , \key_mem[0][111] , \key_mem[0][110] , \key_mem[0][109] , 
       \key_mem[0][108] , \key_mem[0][107] , \key_mem[0][106] , \key_mem[0][105] , 
       \key_mem[0][104] , \key_mem[0][103] , \key_mem[0][102] , \key_mem[0][101] , 
       \key_mem[0][100] , \key_mem[0][99] , \key_mem[0][98] , \key_mem[0][97] , 
       \key_mem[0][96] , \key_mem[0][95] , \key_mem[0][94] , \key_mem[0][93] , 
       \key_mem[0][92] , \key_mem[0][91] , \key_mem[0][90] , \key_mem[0][89] , 
       \key_mem[0][88] , \key_mem[0][87] , \key_mem[0][86] , \key_mem[0][85] , 
       \key_mem[0][84] , \key_mem[0][83] , \key_mem[0][82] , \key_mem[0][81] , 
       \key_mem[0][80] , \key_mem[0][79] , \key_mem[0][78] , \key_mem[0][77] , 
       \key_mem[0][76] , \key_mem[0][75] , \key_mem[0][74] , \key_mem[0][73] , 
       \key_mem[0][72] , \key_mem[0][71] , \key_mem[0][70] , \key_mem[0][69] , 
       \key_mem[0][68] , \key_mem[0][67] , \key_mem[0][66] , \key_mem[0][65] , 
       \key_mem[0][64] , \key_mem[0][63] , \key_mem[0][62] , \key_mem[0][61] , 
       \key_mem[0][60] , \key_mem[0][59] , \key_mem[0][58] , \key_mem[0][57] , 
       \key_mem[0][56] , \key_mem[0][55] , \key_mem[0][54] , \key_mem[0][53] , 
       \key_mem[0][52] , \key_mem[0][51] , \key_mem[0][50] , \key_mem[0][49] , 
       \key_mem[0][48] , \key_mem[0][47] , \key_mem[0][46] , \key_mem[0][45] , 
       \key_mem[0][44] , \key_mem[0][43] , \key_mem[0][42] , \key_mem[0][41] , 
       \key_mem[0][40] , \key_mem[0][39] , \key_mem[0][38] , \key_mem[0][37] , 
       \key_mem[0][36] , \key_mem[0][35] , \key_mem[0][34] , \key_mem[0][33] , 
       \key_mem[0][32] , \key_mem[0][31] , \key_mem[0][30] , \key_mem[0][29] , 
       \key_mem[0][28] , \key_mem[0][27] , \key_mem[0][26] , \key_mem[0][25] , 
       \key_mem[0][24] , \key_mem[0][23] , \key_mem[0][22] , \key_mem[0][21] , 
       \key_mem[0][20] , \key_mem[0][19] , \key_mem[0][18] , \key_mem[0][17] , 
       \key_mem[0][16] , \key_mem[0][15] , \key_mem[0][14] , \key_mem[0][13] , 
       \key_mem[0][12] , \key_mem[0][11] , \key_mem[0][10] , \key_mem[0][9] , 
       \key_mem[0][8] , \key_mem[0][7] , \key_mem[0][6] , \key_mem[0][5] , \key_mem[0][4] 
       , \key_mem[0][3] , \key_mem[0][2] , \key_mem[0][1] , \key_mem[0][0] , 
       \key_mem[1][127] , \key_mem[1][126] , \key_mem[1][125] , \key_mem[1][124] , 
       \key_mem[1][123] , \key_mem[1][122] , \key_mem[1][121] , \key_mem[1][120] , 
       \key_mem[1][119] , \key_mem[1][118] , \key_mem[1][117] , \key_mem[1][116] , 
       \key_mem[1][115] , \key_mem[1][114] , \key_mem[1][113] , \key_mem[1][112] , 
       \key_mem[1][111] , \key_mem[1][110] , \key_mem[1][109] , \key_mem[1][108] , 
       \key_mem[1][107] , \key_mem[1][106] , \key_mem[1][105] , \key_mem[1][104] , 
       \key_mem[1][103] , \key_mem[1][102] , \key_mem[1][101] , \key_mem[1][100] , 
       \key_mem[1][99] , \key_mem[1][98] , \key_mem[1][97] , \key_mem[1][96] , 
       \key_mem[1][95] , \key_mem[1][94] , \key_mem[1][93] , \key_mem[1][92] , 
       \key_mem[1][91] , \key_mem[1][90] , \key_mem[1][89] , \key_mem[1][88] , 
       \key_mem[1][87] , \key_mem[1][86] , \key_mem[1][85] , \key_mem[1][84] , 
       \key_mem[1][83] , \key_mem[1][82] , \key_mem[1][81] , \key_mem[1][80] , 
       \key_mem[1][79] , \key_mem[1][78] , \key_mem[1][77] , \key_mem[1][76] , 
       \key_mem[1][75] , \key_mem[1][74] , \key_mem[1][73] , \key_mem[1][72] , 
       \key_mem[1][71] , \key_mem[1][70] , \key_mem[1][69] , \key_mem[1][68] , 
       \key_mem[1][67] , \key_mem[1][66] , \key_mem[1][65] , \key_mem[1][64] , 
       \key_mem[1][63] , \key_mem[1][62] , \key_mem[1][61] , \key_mem[1][60] , 
       \key_mem[1][59] , \key_mem[1][58] , \key_mem[1][57] , \key_mem[1][56] , 
       \key_mem[1][55] , \key_mem[1][54] , \key_mem[1][53] , \key_mem[1][52] , 
       \key_mem[1][51] , \key_mem[1][50] , \key_mem[1][49] , \key_mem[1][48] , 
       \key_mem[1][47] , \key_mem[1][46] , \key_mem[1][45] , \key_mem[1][44] , 
       \key_mem[1][43] , \key_mem[1][42] , \key_mem[1][41] , \key_mem[1][40] , 
       \key_mem[1][39] , \key_mem[1][38] , \key_mem[1][37] , \key_mem[1][36] , 
       \key_mem[1][35] , \key_mem[1][34] , \key_mem[1][33] , \key_mem[1][32] , 
       \key_mem[1][31] , \key_mem[1][30] , \key_mem[1][29] , \key_mem[1][28] , 
       \key_mem[1][27] , \key_mem[1][26] , \key_mem[1][25] , \key_mem[1][24] , 
       \key_mem[1][23] , \key_mem[1][22] , \key_mem[1][21] , \key_mem[1][20] , 
       \key_mem[1][19] , \key_mem[1][18] , \key_mem[1][17] , \key_mem[1][16] , 
       \key_mem[1][15] , \key_mem[1][14] , \key_mem[1][13] , \key_mem[1][12] , 
       \key_mem[1][11] , \key_mem[1][10] , \key_mem[1][9] , \key_mem[1][8] , 
       \key_mem[1][7] , \key_mem[1][6] , \key_mem[1][5] , \key_mem[1][4] , \key_mem[1][3] 
       , \key_mem[1][2] , \key_mem[1][1] , \key_mem[1][0] , \key_mem[2][127] , 
       \key_mem[2][126] , \key_mem[2][125] , \key_mem[2][124] , \key_mem[2][123] , 
       \key_mem[2][122] , \key_mem[2][121] , \key_mem[2][120] , \key_mem[2][119] , 
       \key_mem[2][118] , \key_mem[2][117] , \key_mem[2][116] , \key_mem[2][115] , 
       \key_mem[2][114] , \key_mem[2][113] , \key_mem[2][112] , \key_mem[2][111] , 
       \key_mem[2][110] , \key_mem[2][109] , \key_mem[2][108] , \key_mem[2][107] , 
       \key_mem[2][106] , \key_mem[2][105] , \key_mem[2][104] , \key_mem[2][103] , 
       \key_mem[2][102] , \key_mem[2][101] , \key_mem[2][100] , \key_mem[2][99] , 
       \key_mem[2][98] , \key_mem[2][97] , \key_mem[2][96] , \key_mem[2][95] , 
       \key_mem[2][94] , \key_mem[2][93] , \key_mem[2][92] , \key_mem[2][91] , 
       \key_mem[2][90] , \key_mem[2][89] , \key_mem[2][88] , \key_mem[2][87] , 
       \key_mem[2][86] , \key_mem[2][85] , \key_mem[2][84] , \key_mem[2][83] , 
       \key_mem[2][82] , \key_mem[2][81] , \key_mem[2][80] , \key_mem[2][79] , 
       \key_mem[2][78] , \key_mem[2][77] , \key_mem[2][76] , \key_mem[2][75] , 
       \key_mem[2][74] , \key_mem[2][73] , \key_mem[2][72] , \key_mem[2][71] , 
       \key_mem[2][70] , \key_mem[2][69] , \key_mem[2][68] , \key_mem[2][67] , 
       \key_mem[2][66] , \key_mem[2][65] , \key_mem[2][64] , \key_mem[2][63] , 
       \key_mem[2][62] , \key_mem[2][61] , \key_mem[2][60] , \key_mem[2][59] , 
       \key_mem[2][58] , \key_mem[2][57] , \key_mem[2][56] , \key_mem[2][55] , 
       \key_mem[2][54] , \key_mem[2][53] , \key_mem[2][52] , \key_mem[2][51] , 
       \key_mem[2][50] , \key_mem[2][49] , \key_mem[2][48] , \key_mem[2][47] , 
       \key_mem[2][46] , \key_mem[2][45] , \key_mem[2][44] , \key_mem[2][43] , 
       \key_mem[2][42] , \key_mem[2][41] , \key_mem[2][40] , \key_mem[2][39] , 
       \key_mem[2][38] , \key_mem[2][37] , \key_mem[2][36] , \key_mem[2][35] , 
       \key_mem[2][34] , \key_mem[2][33] , \key_mem[2][32] , \key_mem[2][31] , 
       \key_mem[2][30] , \key_mem[2][29] , \key_mem[2][28] , \key_mem[2][27] , 
       \key_mem[2][26] , \key_mem[2][25] , \key_mem[2][24] , \key_mem[2][23] , 
       \key_mem[2][22] , \key_mem[2][21] , \key_mem[2][20] , \key_mem[2][19] , 
       \key_mem[2][18] , \key_mem[2][17] , \key_mem[2][16] , \key_mem[2][15] , 
       \key_mem[2][14] , \key_mem[2][13] , \key_mem[2][12] , \key_mem[2][11] , 
       \key_mem[2][10] , \key_mem[2][9] , \key_mem[2][8] , \key_mem[2][7] , 
       \key_mem[2][6] , \key_mem[2][5] , \key_mem[2][4] , \key_mem[2][3] , \key_mem[2][2] 
       , \key_mem[2][1] , \key_mem[2][0] , \key_mem[3][127] , \key_mem[3][126] , 
       \key_mem[3][125] , \key_mem[3][124] , \key_mem[3][123] , \key_mem[3][122] , 
       \key_mem[3][121] , \key_mem[3][120] , \key_mem[3][119] , \key_mem[3][118] , 
       \key_mem[3][117] , \key_mem[3][116] , \key_mem[3][115] , \key_mem[3][114] , 
       \key_mem[3][113] , \key_mem[3][112] , \key_mem[3][111] , \key_mem[3][110] , 
       \key_mem[3][109] , \key_mem[3][108] , \key_mem[3][107] , \key_mem[3][106] , 
       \key_mem[3][105] , \key_mem[3][104] , \key_mem[3][103] , \key_mem[3][102] , 
       \key_mem[3][101] , \key_mem[3][100] , \key_mem[3][99] , \key_mem[3][98] , 
       \key_mem[3][97] , \key_mem[3][96] , \key_mem[3][95] , \key_mem[3][94] , 
       \key_mem[3][93] , \key_mem[3][92] , \key_mem[3][91] , \key_mem[3][90] , 
       \key_mem[3][89] , \key_mem[3][88] , \key_mem[3][87] , \key_mem[3][86] , 
       \key_mem[3][85] , \key_mem[3][84] , \key_mem[3][83] , \key_mem[3][82] , 
       \key_mem[3][81] , \key_mem[3][80] , \key_mem[3][79] , \key_mem[3][78] , 
       \key_mem[3][77] , \key_mem[3][76] , \key_mem[3][75] , \key_mem[3][74] , 
       \key_mem[3][73] , \key_mem[3][72] , \key_mem[3][71] , \key_mem[3][70] , 
       \key_mem[3][69] , \key_mem[3][68] , \key_mem[3][67] , \key_mem[3][66] , 
       \key_mem[3][65] , \key_mem[3][64] , \key_mem[3][63] , \key_mem[3][62] , 
       \key_mem[3][61] , \key_mem[3][60] , \key_mem[3][59] , \key_mem[3][58] , 
       \key_mem[3][57] , \key_mem[3][56] , \key_mem[3][55] , \key_mem[3][54] , 
       \key_mem[3][53] , \key_mem[3][52] , \key_mem[3][51] , \key_mem[3][50] , 
       \key_mem[3][49] , \key_mem[3][48] , \key_mem[3][47] , \key_mem[3][46] , 
       \key_mem[3][45] , \key_mem[3][44] , \key_mem[3][43] , \key_mem[3][42] , 
       \key_mem[3][41] , \key_mem[3][40] , \key_mem[3][39] , \key_mem[3][38] , 
       \key_mem[3][37] , \key_mem[3][36] , \key_mem[3][35] , \key_mem[3][34] , 
       \key_mem[3][33] , \key_mem[3][32] , \key_mem[3][31] , \key_mem[3][30] , 
       \key_mem[3][29] , \key_mem[3][28] , \key_mem[3][27] , \key_mem[3][26] , 
       \key_mem[3][25] , \key_mem[3][24] , \key_mem[3][23] , \key_mem[3][22] , 
       \key_mem[3][21] , \key_mem[3][20] , \key_mem[3][19] , \key_mem[3][18] , 
       \key_mem[3][17] , \key_mem[3][16] , \key_mem[3][15] , \key_mem[3][14] , 
       \key_mem[3][13] , \key_mem[3][12] , \key_mem[3][11] , \key_mem[3][10] , 
       \key_mem[3][9] , \key_mem[3][8] , \key_mem[3][7] , \key_mem[3][6] , \key_mem[3][5] 
       , \key_mem[3][4] , \key_mem[3][3] , \key_mem[3][2] , \key_mem[3][1] , 
       \key_mem[3][0] , \key_mem[4][127] , \key_mem[4][126] , \key_mem[4][125] , 
       \key_mem[4][124] , \key_mem[4][123] , \key_mem[4][122] , \key_mem[4][121] , 
       \key_mem[4][120] , \key_mem[4][119] , \key_mem[4][118] , \key_mem[4][117] , 
       \key_mem[4][116] , \key_mem[4][115] , \key_mem[4][114] , \key_mem[4][113] , 
       \key_mem[4][112] , \key_mem[4][111] , \key_mem[4][110] , \key_mem[4][109] , 
       \key_mem[4][108] , \key_mem[4][107] , \key_mem[4][106] , \key_mem[4][105] , 
       \key_mem[4][104] , \key_mem[4][103] , \key_mem[4][102] , \key_mem[4][101] , 
       \key_mem[4][100] , \key_mem[4][99] , \key_mem[4][98] , \key_mem[4][97] , 
       \key_mem[4][96] , \key_mem[4][95] , \key_mem[4][94] , \key_mem[4][93] , 
       \key_mem[4][92] , \key_mem[4][91] , \key_mem[4][90] , \key_mem[4][89] , 
       \key_mem[4][88] , \key_mem[4][87] , \key_mem[4][86] , \key_mem[4][85] , 
       \key_mem[4][84] , \key_mem[4][83] , \key_mem[4][82] , \key_mem[4][81] , 
       \key_mem[4][80] , \key_mem[4][79] , \key_mem[4][78] , \key_mem[4][77] , 
       \key_mem[4][76] , \key_mem[4][75] , \key_mem[4][74] , \key_mem[4][73] , 
       \key_mem[4][72] , \key_mem[4][71] , \key_mem[4][70] , \key_mem[4][69] , 
       \key_mem[4][68] , \key_mem[4][67] , \key_mem[4][66] , \key_mem[4][65] , 
       \key_mem[4][64] , \key_mem[4][63] , \key_mem[4][62] , \key_mem[4][61] , 
       \key_mem[4][60] , \key_mem[4][59] , \key_mem[4][58] , \key_mem[4][57] , 
       \key_mem[4][56] , \key_mem[4][55] , \key_mem[4][54] , \key_mem[4][53] , 
       \key_mem[4][52] , \key_mem[4][51] , \key_mem[4][50] , \key_mem[4][49] , 
       \key_mem[4][48] , \key_mem[4][47] , \key_mem[4][46] , \key_mem[4][45] , 
       \key_mem[4][44] , \key_mem[4][43] , \key_mem[4][42] , \key_mem[4][41] , 
       \key_mem[4][40] , \key_mem[4][39] , \key_mem[4][38] , \key_mem[4][37] , 
       \key_mem[4][36] , \key_mem[4][35] , \key_mem[4][34] , \key_mem[4][33] , 
       \key_mem[4][32] , \key_mem[4][31] , \key_mem[4][30] , \key_mem[4][29] , 
       \key_mem[4][28] , \key_mem[4][27] , \key_mem[4][26] , \key_mem[4][25] , 
       \key_mem[4][24] , \key_mem[4][23] , \key_mem[4][22] , \key_mem[4][21] , 
       \key_mem[4][20] , \key_mem[4][19] , \key_mem[4][18] , \key_mem[4][17] , 
       \key_mem[4][16] , \key_mem[4][15] , \key_mem[4][14] , \key_mem[4][13] , 
       \key_mem[4][12] , \key_mem[4][11] , \key_mem[4][10] , \key_mem[4][9] , 
       \key_mem[4][8] , \key_mem[4][7] , \key_mem[4][6] , \key_mem[4][5] , \key_mem[4][4] 
       , \key_mem[4][3] , \key_mem[4][2] , \key_mem[4][1] , \key_mem[4][0] , 
       \key_mem[5][127] , \key_mem[5][126] , \key_mem[5][125] , \key_mem[5][124] , 
       \key_mem[5][123] , \key_mem[5][122] , \key_mem[5][121] , \key_mem[5][120] , 
       \key_mem[5][119] , \key_mem[5][118] , \key_mem[5][117] , \key_mem[5][116] , 
       \key_mem[5][115] , \key_mem[5][114] , \key_mem[5][113] , \key_mem[5][112] , 
       \key_mem[5][111] , \key_mem[5][110] , \key_mem[5][109] , \key_mem[5][108] , 
       \key_mem[5][107] , \key_mem[5][106] , \key_mem[5][105] , \key_mem[5][104] , 
       \key_mem[5][103] , \key_mem[5][102] , \key_mem[5][101] , \key_mem[5][100] , 
       \key_mem[5][99] , \key_mem[5][98] , \key_mem[5][97] , \key_mem[5][96] , 
       \key_mem[5][95] , \key_mem[5][94] , \key_mem[5][93] , \key_mem[5][92] , 
       \key_mem[5][91] , \key_mem[5][90] , \key_mem[5][89] , \key_mem[5][88] , 
       \key_mem[5][87] , \key_mem[5][86] , \key_mem[5][85] , \key_mem[5][84] , 
       \key_mem[5][83] , \key_mem[5][82] , \key_mem[5][81] , \key_mem[5][80] , 
       \key_mem[5][79] , \key_mem[5][78] , \key_mem[5][77] , \key_mem[5][76] , 
       \key_mem[5][75] , \key_mem[5][74] , \key_mem[5][73] , \key_mem[5][72] , 
       \key_mem[5][71] , \key_mem[5][70] , \key_mem[5][69] , \key_mem[5][68] , 
       \key_mem[5][67] , \key_mem[5][66] , \key_mem[5][65] , \key_mem[5][64] , 
       \key_mem[5][63] , \key_mem[5][62] , \key_mem[5][61] , \key_mem[5][60] , 
       \key_mem[5][59] , \key_mem[5][58] , \key_mem[5][57] , \key_mem[5][56] , 
       \key_mem[5][55] , \key_mem[5][54] , \key_mem[5][53] , \key_mem[5][52] , 
       \key_mem[5][51] , \key_mem[5][50] , \key_mem[5][49] , \key_mem[5][48] , 
       \key_mem[5][47] , \key_mem[5][46] , \key_mem[5][45] , \key_mem[5][44] , 
       \key_mem[5][43] , \key_mem[5][42] , \key_mem[5][41] , \key_mem[5][40] , 
       \key_mem[5][39] , \key_mem[5][38] , \key_mem[5][37] , \key_mem[5][36] , 
       \key_mem[5][35] , \key_mem[5][34] , \key_mem[5][33] , \key_mem[5][32] , 
       \key_mem[5][31] , \key_mem[5][30] , \key_mem[5][29] , \key_mem[5][28] , 
       \key_mem[5][27] , \key_mem[5][26] , \key_mem[5][25] , \key_mem[5][24] , 
       \key_mem[5][23] , \key_mem[5][22] , \key_mem[5][21] , \key_mem[5][20] , 
       \key_mem[5][19] , \key_mem[5][18] , \key_mem[5][17] , \key_mem[5][16] , 
       \key_mem[5][15] , \key_mem[5][14] , \key_mem[5][13] , \key_mem[5][12] , 
       \key_mem[5][11] , \key_mem[5][10] , \key_mem[5][9] , \key_mem[5][8] , 
       \key_mem[5][7] , \key_mem[5][6] , \key_mem[5][5] , \key_mem[5][4] , \key_mem[5][3] 
       , \key_mem[5][2] , \key_mem[5][1] , \key_mem[5][0] , \key_mem[6][127] , 
       \key_mem[6][126] , \key_mem[6][125] , \key_mem[6][124] , \key_mem[6][123] , 
       \key_mem[6][122] , \key_mem[6][121] , \key_mem[6][120] , \key_mem[6][119] , 
       \key_mem[6][118] , \key_mem[6][117] , \key_mem[6][116] , \key_mem[6][115] , 
       \key_mem[6][114] , \key_mem[6][113] , \key_mem[6][112] , \key_mem[6][111] , 
       \key_mem[6][110] , \key_mem[6][109] , \key_mem[6][108] , \key_mem[6][107] , 
       \key_mem[6][106] , \key_mem[6][105] , \key_mem[6][104] , \key_mem[6][103] , 
       \key_mem[6][102] , \key_mem[6][101] , \key_mem[6][100] , \key_mem[6][99] , 
       \key_mem[6][98] , \key_mem[6][97] , \key_mem[6][96] , \key_mem[6][95] , 
       \key_mem[6][94] , \key_mem[6][93] , \key_mem[6][92] , \key_mem[6][91] , 
       \key_mem[6][90] , \key_mem[6][89] , \key_mem[6][88] , \key_mem[6][87] , 
       \key_mem[6][86] , \key_mem[6][85] , \key_mem[6][84] , \key_mem[6][83] , 
       \key_mem[6][82] , \key_mem[6][81] , \key_mem[6][80] , \key_mem[6][79] , 
       \key_mem[6][78] , \key_mem[6][77] , \key_mem[6][76] , \key_mem[6][75] , 
       \key_mem[6][74] , \key_mem[6][73] , \key_mem[6][72] , \key_mem[6][71] , 
       \key_mem[6][70] , \key_mem[6][69] , \key_mem[6][68] , \key_mem[6][67] , 
       \key_mem[6][66] , \key_mem[6][65] , \key_mem[6][64] , \key_mem[6][63] , 
       \key_mem[6][62] , \key_mem[6][61] , \key_mem[6][60] , \key_mem[6][59] , 
       \key_mem[6][58] , \key_mem[6][57] , \key_mem[6][56] , \key_mem[6][55] , 
       \key_mem[6][54] , \key_mem[6][53] , \key_mem[6][52] , \key_mem[6][51] , 
       \key_mem[6][50] , \key_mem[6][49] , \key_mem[6][48] , \key_mem[6][47] , 
       \key_mem[6][46] , \key_mem[6][45] , \key_mem[6][44] , \key_mem[6][43] , 
       \key_mem[6][42] , \key_mem[6][41] , \key_mem[6][40] , \key_mem[6][39] , 
       \key_mem[6][38] , \key_mem[6][37] , \key_mem[6][36] , \key_mem[6][35] , 
       \key_mem[6][34] , \key_mem[6][33] , \key_mem[6][32] , \key_mem[6][31] , 
       \key_mem[6][30] , \key_mem[6][29] , \key_mem[6][28] , \key_mem[6][27] , 
       \key_mem[6][26] , \key_mem[6][25] , \key_mem[6][24] , \key_mem[6][23] , 
       \key_mem[6][22] , \key_mem[6][21] , \key_mem[6][20] , \key_mem[6][19] , 
       \key_mem[6][18] , \key_mem[6][17] , \key_mem[6][16] , \key_mem[6][15] , 
       \key_mem[6][14] , \key_mem[6][13] , \key_mem[6][12] , \key_mem[6][11] , 
       \key_mem[6][10] , \key_mem[6][9] , \key_mem[6][8] , \key_mem[6][7] , 
       \key_mem[6][6] , \key_mem[6][5] , \key_mem[6][4] , \key_mem[6][3] , \key_mem[6][2] 
       , \key_mem[6][1] , \key_mem[6][0] , \key_mem[7][127] , \key_mem[7][126] , 
       \key_mem[7][125] , \key_mem[7][124] , \key_mem[7][123] , \key_mem[7][122] , 
       \key_mem[7][121] , \key_mem[7][120] , \key_mem[7][119] , \key_mem[7][118] , 
       \key_mem[7][117] , \key_mem[7][116] , \key_mem[7][115] , \key_mem[7][114] , 
       \key_mem[7][113] , \key_mem[7][112] , \key_mem[7][111] , \key_mem[7][110] , 
       \key_mem[7][109] , \key_mem[7][108] , \key_mem[7][107] , \key_mem[7][106] , 
       \key_mem[7][105] , \key_mem[7][104] , \key_mem[7][103] , \key_mem[7][102] , 
       \key_mem[7][101] , \key_mem[7][100] , \key_mem[7][99] , \key_mem[7][98] , 
       \key_mem[7][97] , \key_mem[7][96] , \key_mem[7][95] , \key_mem[7][94] , 
       \key_mem[7][93] , \key_mem[7][92] , \key_mem[7][91] , \key_mem[7][90] , 
       \key_mem[7][89] , \key_mem[7][88] , \key_mem[7][87] , \key_mem[7][86] , 
       \key_mem[7][85] , \key_mem[7][84] , \key_mem[7][83] , \key_mem[7][82] , 
       \key_mem[7][81] , \key_mem[7][80] , \key_mem[7][79] , \key_mem[7][78] , 
       \key_mem[7][77] , \key_mem[7][76] , \key_mem[7][75] , \key_mem[7][74] , 
       \key_mem[7][73] , \key_mem[7][72] , \key_mem[7][71] , \key_mem[7][70] , 
       \key_mem[7][69] , \key_mem[7][68] , \key_mem[7][67] , \key_mem[7][66] , 
       \key_mem[7][65] , \key_mem[7][64] , \key_mem[7][63] , \key_mem[7][62] , 
       \key_mem[7][61] , \key_mem[7][60] , \key_mem[7][59] , \key_mem[7][58] , 
       \key_mem[7][57] , \key_mem[7][56] , \key_mem[7][55] , \key_mem[7][54] , 
       \key_mem[7][53] , \key_mem[7][52] , \key_mem[7][51] , \key_mem[7][50] , 
       \key_mem[7][49] , \key_mem[7][48] , \key_mem[7][47] , \key_mem[7][46] , 
       \key_mem[7][45] , \key_mem[7][44] , \key_mem[7][43] , \key_mem[7][42] , 
       \key_mem[7][41] , \key_mem[7][40] , \key_mem[7][39] , \key_mem[7][38] , 
       \key_mem[7][37] , \key_mem[7][36] , \key_mem[7][35] , \key_mem[7][34] , 
       \key_mem[7][33] , \key_mem[7][32] , \key_mem[7][31] , \key_mem[7][30] , 
       \key_mem[7][29] , \key_mem[7][28] , \key_mem[7][27] , \key_mem[7][26] , 
       \key_mem[7][25] , \key_mem[7][24] , \key_mem[7][23] , \key_mem[7][22] , 
       \key_mem[7][21] , \key_mem[7][20] , \key_mem[7][19] , \key_mem[7][18] , 
       \key_mem[7][17] , \key_mem[7][16] , \key_mem[7][15] , \key_mem[7][14] , 
       \key_mem[7][13] , \key_mem[7][12] , \key_mem[7][11] , \key_mem[7][10] , 
       \key_mem[7][9] , \key_mem[7][8] , \key_mem[7][7] , \key_mem[7][6] , \key_mem[7][5] 
       , \key_mem[7][4] , \key_mem[7][3] , \key_mem[7][2] , \key_mem[7][1] , 
       \key_mem[7][0] , \key_mem[8][127] , \key_mem[8][126] , \key_mem[8][125] , 
       \key_mem[8][124] , \key_mem[8][123] , \key_mem[8][122] , \key_mem[8][121] , 
       \key_mem[8][120] , \key_mem[8][119] , \key_mem[8][118] , \key_mem[8][117] , 
       \key_mem[8][116] , \key_mem[8][115] , \key_mem[8][114] , \key_mem[8][113] , 
       \key_mem[8][112] , \key_mem[8][111] , \key_mem[8][110] , \key_mem[8][109] , 
       \key_mem[8][108] , \key_mem[8][107] , \key_mem[8][106] , \key_mem[8][105] , 
       \key_mem[8][104] , \key_mem[8][103] , \key_mem[8][102] , \key_mem[8][101] , 
       \key_mem[8][100] , \key_mem[8][99] , \key_mem[8][98] , \key_mem[8][97] , 
       \key_mem[8][96] , \key_mem[8][95] , \key_mem[8][94] , \key_mem[8][93] , 
       \key_mem[8][92] , \key_mem[8][91] , \key_mem[8][90] , \key_mem[8][89] , 
       \key_mem[8][88] , \key_mem[8][87] , \key_mem[8][86] , \key_mem[8][85] , 
       \key_mem[8][84] , \key_mem[8][83] , \key_mem[8][82] , \key_mem[8][81] , 
       \key_mem[8][80] , \key_mem[8][79] , \key_mem[8][78] , \key_mem[8][77] , 
       \key_mem[8][76] , \key_mem[8][75] , \key_mem[8][74] , \key_mem[8][73] , 
       \key_mem[8][72] , \key_mem[8][71] , \key_mem[8][70] , \key_mem[8][69] , 
       \key_mem[8][68] , \key_mem[8][67] , \key_mem[8][66] , \key_mem[8][65] , 
       \key_mem[8][64] , \key_mem[8][63] , \key_mem[8][62] , \key_mem[8][61] , 
       \key_mem[8][60] , \key_mem[8][59] , \key_mem[8][58] , \key_mem[8][57] , 
       \key_mem[8][56] , \key_mem[8][55] , \key_mem[8][54] , \key_mem[8][53] , 
       \key_mem[8][52] , \key_mem[8][51] , \key_mem[8][50] , \key_mem[8][49] , 
       \key_mem[8][48] , \key_mem[8][47] , \key_mem[8][46] , \key_mem[8][45] , 
       \key_mem[8][44] , \key_mem[8][43] , \key_mem[8][42] , \key_mem[8][41] , 
       \key_mem[8][40] , \key_mem[8][39] , \key_mem[8][38] , \key_mem[8][37] , 
       \key_mem[8][36] , \key_mem[8][35] , \key_mem[8][34] , \key_mem[8][33] , 
       \key_mem[8][32] , \key_mem[8][31] , \key_mem[8][30] , \key_mem[8][29] , 
       \key_mem[8][28] , \key_mem[8][27] , \key_mem[8][26] , \key_mem[8][25] , 
       \key_mem[8][24] , \key_mem[8][23] , \key_mem[8][22] , \key_mem[8][21] , 
       \key_mem[8][20] , \key_mem[8][19] , \key_mem[8][18] , \key_mem[8][17] , 
       \key_mem[8][16] , \key_mem[8][15] , \key_mem[8][14] , \key_mem[8][13] , 
       \key_mem[8][12] , \key_mem[8][11] , \key_mem[8][10] , \key_mem[8][9] , 
       \key_mem[8][8] , \key_mem[8][7] , \key_mem[8][6] , \key_mem[8][5] , \key_mem[8][4] 
       , \key_mem[8][3] , \key_mem[8][2] , \key_mem[8][1] , \key_mem[8][0] , 
       \key_mem[9][127] , \key_mem[9][126] , \key_mem[9][125] , \key_mem[9][124] , 
       \key_mem[9][123] , \key_mem[9][122] , \key_mem[9][121] , \key_mem[9][120] , 
       \key_mem[9][119] , \key_mem[9][118] , \key_mem[9][117] , \key_mem[9][116] , 
       \key_mem[9][115] , \key_mem[9][114] , \key_mem[9][113] , \key_mem[9][112] , 
       \key_mem[9][111] , \key_mem[9][110] , \key_mem[9][109] , \key_mem[9][108] , 
       \key_mem[9][107] , \key_mem[9][106] , \key_mem[9][105] , \key_mem[9][104] , 
       \key_mem[9][103] , \key_mem[9][102] , \key_mem[9][101] , \key_mem[9][100] , 
       \key_mem[9][99] , \key_mem[9][98] , \key_mem[9][97] , \key_mem[9][96] , 
       \key_mem[9][95] , \key_mem[9][94] , \key_mem[9][93] , \key_mem[9][92] , 
       \key_mem[9][91] , \key_mem[9][90] , \key_mem[9][89] , \key_mem[9][88] , 
       \key_mem[9][87] , \key_mem[9][86] , \key_mem[9][85] , \key_mem[9][84] , 
       \key_mem[9][83] , \key_mem[9][82] , \key_mem[9][81] , \key_mem[9][80] , 
       \key_mem[9][79] , \key_mem[9][78] , \key_mem[9][77] , \key_mem[9][76] , 
       \key_mem[9][75] , \key_mem[9][74] , \key_mem[9][73] , \key_mem[9][72] , 
       \key_mem[9][71] , \key_mem[9][70] , \key_mem[9][69] , \key_mem[9][68] , 
       \key_mem[9][67] , \key_mem[9][66] , \key_mem[9][65] , \key_mem[9][64] , 
       \key_mem[9][63] , \key_mem[9][62] , \key_mem[9][61] , \key_mem[9][60] , 
       \key_mem[9][59] , \key_mem[9][58] , \key_mem[9][57] , \key_mem[9][56] , 
       \key_mem[9][55] , \key_mem[9][54] , \key_mem[9][53] , \key_mem[9][52] , 
       \key_mem[9][51] , \key_mem[9][50] , \key_mem[9][49] , \key_mem[9][48] , 
       \key_mem[9][47] , \key_mem[9][46] , \key_mem[9][45] , \key_mem[9][44] , 
       \key_mem[9][43] , \key_mem[9][42] , \key_mem[9][41] , \key_mem[9][40] , 
       \key_mem[9][39] , \key_mem[9][38] , \key_mem[9][37] , \key_mem[9][36] , 
       \key_mem[9][35] , \key_mem[9][34] , \key_mem[9][33] , \key_mem[9][32] , 
       \key_mem[9][31] , \key_mem[9][30] , \key_mem[9][29] , \key_mem[9][28] , 
       \key_mem[9][27] , \key_mem[9][26] , \key_mem[9][25] , \key_mem[9][24] , 
       \key_mem[9][23] , \key_mem[9][22] , \key_mem[9][21] , \key_mem[9][20] , 
       \key_mem[9][19] , \key_mem[9][18] , \key_mem[9][17] , \key_mem[9][16] , 
       \key_mem[9][15] , \key_mem[9][14] , \key_mem[9][13] , \key_mem[9][12] , 
       \key_mem[9][11] , \key_mem[9][10] , \key_mem[9][9] , \key_mem[9][8] , 
       \key_mem[9][7] , \key_mem[9][6] , \key_mem[9][5] , \key_mem[9][4] , \key_mem[9][3] 
       , \key_mem[9][2] , \key_mem[9][1] , \key_mem[9][0] , \key_mem[10][127] , 
       \key_mem[10][126] , \key_mem[10][125] , \key_mem[10][124] , \key_mem[10][123] , 
       \key_mem[10][122] , \key_mem[10][121] , \key_mem[10][120] , \key_mem[10][119] , 
       \key_mem[10][118] , \key_mem[10][117] , \key_mem[10][116] , \key_mem[10][115] , 
       \key_mem[10][114] , \key_mem[10][113] , \key_mem[10][112] , \key_mem[10][111] , 
       \key_mem[10][110] , \key_mem[10][109] , \key_mem[10][108] , \key_mem[10][107] , 
       \key_mem[10][106] , \key_mem[10][105] , \key_mem[10][104] , \key_mem[10][103] , 
       \key_mem[10][102] , \key_mem[10][101] , \key_mem[10][100] , \key_mem[10][99] , 
       \key_mem[10][98] , \key_mem[10][97] , \key_mem[10][96] , \key_mem[10][95] , 
       \key_mem[10][94] , \key_mem[10][93] , \key_mem[10][92] , \key_mem[10][91] , 
       \key_mem[10][90] , \key_mem[10][89] , \key_mem[10][88] , \key_mem[10][87] , 
       \key_mem[10][86] , \key_mem[10][85] , \key_mem[10][84] , \key_mem[10][83] , 
       \key_mem[10][82] , \key_mem[10][81] , \key_mem[10][80] , \key_mem[10][79] , 
       \key_mem[10][78] , \key_mem[10][77] , \key_mem[10][76] , \key_mem[10][75] , 
       \key_mem[10][74] , \key_mem[10][73] , \key_mem[10][72] , \key_mem[10][71] , 
       \key_mem[10][70] , \key_mem[10][69] , \key_mem[10][68] , \key_mem[10][67] , 
       \key_mem[10][66] , \key_mem[10][65] , \key_mem[10][64] , \key_mem[10][63] , 
       \key_mem[10][62] , \key_mem[10][61] , \key_mem[10][60] , \key_mem[10][59] , 
       \key_mem[10][58] , \key_mem[10][57] , \key_mem[10][56] , \key_mem[10][55] , 
       \key_mem[10][54] , \key_mem[10][53] , \key_mem[10][52] , \key_mem[10][51] , 
       \key_mem[10][50] , \key_mem[10][49] , \key_mem[10][48] , \key_mem[10][47] , 
       \key_mem[10][46] , \key_mem[10][45] , \key_mem[10][44] , \key_mem[10][43] , 
       \key_mem[10][42] , \key_mem[10][41] , \key_mem[10][40] , \key_mem[10][39] , 
       \key_mem[10][38] , \key_mem[10][37] , \key_mem[10][36] , \key_mem[10][35] , 
       \key_mem[10][34] , \key_mem[10][33] , \key_mem[10][32] , \key_mem[10][31] , 
       \key_mem[10][30] , \key_mem[10][29] , \key_mem[10][28] , \key_mem[10][27] , 
       \key_mem[10][26] , \key_mem[10][25] , \key_mem[10][24] , \key_mem[10][23] , 
       \key_mem[10][22] , \key_mem[10][21] , \key_mem[10][20] , \key_mem[10][19] , 
       \key_mem[10][18] , \key_mem[10][17] , \key_mem[10][16] , \key_mem[10][15] , 
       \key_mem[10][14] , \key_mem[10][13] , \key_mem[10][12] , \key_mem[10][11] , 
       \key_mem[10][10] , \key_mem[10][9] , \key_mem[10][8] , \key_mem[10][7] , 
       \key_mem[10][6] , \key_mem[10][5] , \key_mem[10][4] , \key_mem[10][3] , 
       \key_mem[10][2] , \key_mem[10][1] , \key_mem[10][0] , \key_mem[11][127] , 
       \key_mem[11][126] , \key_mem[11][125] , \key_mem[11][124] , \key_mem[11][123] , 
       \key_mem[11][122] , \key_mem[11][121] , \key_mem[11][120] , \key_mem[11][119] , 
       \key_mem[11][118] , \key_mem[11][117] , \key_mem[11][116] , \key_mem[11][115] , 
       \key_mem[11][114] , \key_mem[11][113] , \key_mem[11][112] , \key_mem[11][111] , 
       \key_mem[11][110] , \key_mem[11][109] , \key_mem[11][108] , \key_mem[11][107] , 
       \key_mem[11][106] , \key_mem[11][105] , \key_mem[11][104] , \key_mem[11][103] , 
       \key_mem[11][102] , \key_mem[11][101] , \key_mem[11][100] , \key_mem[11][99] , 
       \key_mem[11][98] , \key_mem[11][97] , \key_mem[11][96] , \key_mem[11][95] , 
       \key_mem[11][94] , \key_mem[11][93] , \key_mem[11][92] , \key_mem[11][91] , 
       \key_mem[11][90] , \key_mem[11][89] , \key_mem[11][88] , \key_mem[11][87] , 
       \key_mem[11][86] , \key_mem[11][85] , \key_mem[11][84] , \key_mem[11][83] , 
       \key_mem[11][82] , \key_mem[11][81] , \key_mem[11][80] , \key_mem[11][79] , 
       \key_mem[11][78] , \key_mem[11][77] , \key_mem[11][76] , \key_mem[11][75] , 
       \key_mem[11][74] , \key_mem[11][73] , \key_mem[11][72] , \key_mem[11][71] , 
       \key_mem[11][70] , \key_mem[11][69] , \key_mem[11][68] , \key_mem[11][67] , 
       \key_mem[11][66] , \key_mem[11][65] , \key_mem[11][64] , \key_mem[11][63] , 
       \key_mem[11][62] , \key_mem[11][61] , \key_mem[11][60] , \key_mem[11][59] , 
       \key_mem[11][58] , \key_mem[11][57] , \key_mem[11][56] , \key_mem[11][55] , 
       \key_mem[11][54] , \key_mem[11][53] , \key_mem[11][52] , \key_mem[11][51] , 
       \key_mem[11][50] , \key_mem[11][49] , \key_mem[11][48] , \key_mem[11][47] , 
       \key_mem[11][46] , \key_mem[11][45] , \key_mem[11][44] , \key_mem[11][43] , 
       \key_mem[11][42] , \key_mem[11][41] , \key_mem[11][40] , \key_mem[11][39] , 
       \key_mem[11][38] , \key_mem[11][37] , \key_mem[11][36] , \key_mem[11][35] , 
       \key_mem[11][34] , \key_mem[11][33] , \key_mem[11][32] , \key_mem[11][31] , 
       \key_mem[11][30] , \key_mem[11][29] , \key_mem[11][28] , \key_mem[11][27] , 
       \key_mem[11][26] , \key_mem[11][25] , \key_mem[11][24] , \key_mem[11][23] , 
       \key_mem[11][22] , \key_mem[11][21] , \key_mem[11][20] , \key_mem[11][19] , 
       \key_mem[11][18] , \key_mem[11][17] , \key_mem[11][16] , \key_mem[11][15] , 
       \key_mem[11][14] , \key_mem[11][13] , \key_mem[11][12] , \key_mem[11][11] , 
       \key_mem[11][10] , \key_mem[11][9] , \key_mem[11][8] , \key_mem[11][7] , 
       \key_mem[11][6] , \key_mem[11][5] , \key_mem[11][4] , \key_mem[11][3] , 
       \key_mem[11][2] , \key_mem[11][1] , \key_mem[11][0] , \key_mem[12][127] , 
       \key_mem[12][126] , \key_mem[12][125] , \key_mem[12][124] , \key_mem[12][123] , 
       \key_mem[12][122] , \key_mem[12][121] , \key_mem[12][120] , \key_mem[12][119] , 
       \key_mem[12][118] , \key_mem[12][117] , \key_mem[12][116] , \key_mem[12][115] , 
       \key_mem[12][114] , \key_mem[12][113] , \key_mem[12][112] , \key_mem[12][111] , 
       \key_mem[12][110] , \key_mem[12][109] , \key_mem[12][108] , \key_mem[12][107] , 
       \key_mem[12][106] , \key_mem[12][105] , \key_mem[12][104] , \key_mem[12][103] , 
       \key_mem[12][102] , \key_mem[12][101] , \key_mem[12][100] , \key_mem[12][99] , 
       \key_mem[12][98] , \key_mem[12][97] , \key_mem[12][96] , \key_mem[12][95] , 
       \key_mem[12][94] , \key_mem[12][93] , \key_mem[12][92] , \key_mem[12][91] , 
       \key_mem[12][90] , \key_mem[12][89] , \key_mem[12][88] , \key_mem[12][87] , 
       \key_mem[12][86] , \key_mem[12][85] , \key_mem[12][84] , \key_mem[12][83] , 
       \key_mem[12][82] , \key_mem[12][81] , \key_mem[12][80] , \key_mem[12][79] , 
       \key_mem[12][78] , \key_mem[12][77] , \key_mem[12][76] , \key_mem[12][75] , 
       \key_mem[12][74] , \key_mem[12][73] , \key_mem[12][72] , \key_mem[12][71] , 
       \key_mem[12][70] , \key_mem[12][69] , \key_mem[12][68] , \key_mem[12][67] , 
       \key_mem[12][66] , \key_mem[12][65] , \key_mem[12][64] , \key_mem[12][63] , 
       \key_mem[12][62] , \key_mem[12][61] , \key_mem[12][60] , \key_mem[12][59] , 
       \key_mem[12][58] , \key_mem[12][57] , \key_mem[12][56] , \key_mem[12][55] , 
       \key_mem[12][54] , \key_mem[12][53] , \key_mem[12][52] , \key_mem[12][51] , 
       \key_mem[12][50] , \key_mem[12][49] , \key_mem[12][48] , \key_mem[12][47] , 
       \key_mem[12][46] , \key_mem[12][45] , \key_mem[12][44] , \key_mem[12][43] , 
       \key_mem[12][42] , \key_mem[12][41] , \key_mem[12][40] , \key_mem[12][39] , 
       \key_mem[12][38] , \key_mem[12][37] , \key_mem[12][36] , \key_mem[12][35] , 
       \key_mem[12][34] , \key_mem[12][33] , \key_mem[12][32] , \key_mem[12][31] , 
       \key_mem[12][30] , \key_mem[12][29] , \key_mem[12][28] , \key_mem[12][27] , 
       \key_mem[12][26] , \key_mem[12][25] , \key_mem[12][24] , \key_mem[12][23] , 
       \key_mem[12][22] , \key_mem[12][21] , \key_mem[12][20] , \key_mem[12][19] , 
       \key_mem[12][18] , \key_mem[12][17] , \key_mem[12][16] , \key_mem[12][15] , 
       \key_mem[12][14] , \key_mem[12][13] , \key_mem[12][12] , \key_mem[12][11] , 
       \key_mem[12][10] , \key_mem[12][9] , \key_mem[12][8] , \key_mem[12][7] , 
       \key_mem[12][6] , \key_mem[12][5] , \key_mem[12][4] , \key_mem[12][3] , 
       \key_mem[12][2] , \key_mem[12][1] , \key_mem[12][0] , \key_mem[13][127] , 
       \key_mem[13][126] , \key_mem[13][125] , \key_mem[13][124] , \key_mem[13][123] , 
       \key_mem[13][122] , \key_mem[13][121] , \key_mem[13][120] , \key_mem[13][119] , 
       \key_mem[13][118] , \key_mem[13][117] , \key_mem[13][116] , \key_mem[13][115] , 
       \key_mem[13][114] , \key_mem[13][113] , \key_mem[13][112] , \key_mem[13][111] , 
       \key_mem[13][110] , \key_mem[13][109] , \key_mem[13][108] , \key_mem[13][107] , 
       \key_mem[13][106] , \key_mem[13][105] , \key_mem[13][104] , \key_mem[13][103] , 
       \key_mem[13][102] , \key_mem[13][101] , \key_mem[13][100] , \key_mem[13][99] , 
       \key_mem[13][98] , \key_mem[13][97] , \key_mem[13][96] , \key_mem[13][95] , 
       \key_mem[13][94] , \key_mem[13][93] , \key_mem[13][92] , \key_mem[13][91] , 
       \key_mem[13][90] , \key_mem[13][89] , \key_mem[13][88] , \key_mem[13][87] , 
       \key_mem[13][86] , \key_mem[13][85] , \key_mem[13][84] , \key_mem[13][83] , 
       \key_mem[13][82] , \key_mem[13][81] , \key_mem[13][80] , \key_mem[13][79] , 
       \key_mem[13][78] , \key_mem[13][77] , \key_mem[13][76] , \key_mem[13][75] , 
       \key_mem[13][74] , \key_mem[13][73] , \key_mem[13][72] , \key_mem[13][71] , 
       \key_mem[13][70] , \key_mem[13][69] , \key_mem[13][68] , \key_mem[13][67] , 
       \key_mem[13][66] , \key_mem[13][65] , \key_mem[13][64] , \key_mem[13][63] , 
       \key_mem[13][62] , \key_mem[13][61] , \key_mem[13][60] , \key_mem[13][59] , 
       \key_mem[13][58] , \key_mem[13][57] , \key_mem[13][56] , \key_mem[13][55] , 
       \key_mem[13][54] , \key_mem[13][53] , \key_mem[13][52] , \key_mem[13][51] , 
       \key_mem[13][50] , \key_mem[13][49] , \key_mem[13][48] , \key_mem[13][47] , 
       \key_mem[13][46] , \key_mem[13][45] , \key_mem[13][44] , \key_mem[13][43] , 
       \key_mem[13][42] , \key_mem[13][41] , \key_mem[13][40] , \key_mem[13][39] , 
       \key_mem[13][38] , \key_mem[13][37] , \key_mem[13][36] , \key_mem[13][35] , 
       \key_mem[13][34] , \key_mem[13][33] , \key_mem[13][32] , \key_mem[13][31] , 
       \key_mem[13][30] , \key_mem[13][29] , \key_mem[13][28] , \key_mem[13][27] , 
       \key_mem[13][26] , \key_mem[13][25] , \key_mem[13][24] , \key_mem[13][23] , 
       \key_mem[13][22] , \key_mem[13][21] , \key_mem[13][20] , \key_mem[13][19] , 
       \key_mem[13][18] , \key_mem[13][17] , \key_mem[13][16] , \key_mem[13][15] , 
       \key_mem[13][14] , \key_mem[13][13] , \key_mem[13][12] , \key_mem[13][11] , 
       \key_mem[13][10] , \key_mem[13][9] , \key_mem[13][8] , \key_mem[13][7] , 
       \key_mem[13][6] , \key_mem[13][5] , \key_mem[13][4] , \key_mem[13][3] , 
       \key_mem[13][2] , \key_mem[13][1] , \key_mem[13][0] , \key_mem[14][127] , 
       \key_mem[14][126] , \key_mem[14][125] , \key_mem[14][124] , \key_mem[14][123] , 
       \key_mem[14][122] , \key_mem[14][121] , \key_mem[14][120] , \key_mem[14][119] , 
       \key_mem[14][118] , \key_mem[14][117] , \key_mem[14][116] , \key_mem[14][115] , 
       \key_mem[14][114] , \key_mem[14][113] , \key_mem[14][112] , \key_mem[14][111] , 
       \key_mem[14][110] , \key_mem[14][109] , \key_mem[14][108] , \key_mem[14][107] , 
       \key_mem[14][106] , \key_mem[14][105] , \key_mem[14][104] , \key_mem[14][103] , 
       \key_mem[14][102] , \key_mem[14][101] , \key_mem[14][100] , \key_mem[14][99] , 
       \key_mem[14][98] , \key_mem[14][97] , \key_mem[14][96] , \key_mem[14][95] , 
       \key_mem[14][94] , \key_mem[14][93] , \key_mem[14][92] , \key_mem[14][91] , 
       \key_mem[14][90] , \key_mem[14][89] , \key_mem[14][88] , \key_mem[14][87] , 
       \key_mem[14][86] , \key_mem[14][85] , \key_mem[14][84] , \key_mem[14][83] , 
       \key_mem[14][82] , \key_mem[14][81] , \key_mem[14][80] , \key_mem[14][79] , 
       \key_mem[14][78] , \key_mem[14][77] , \key_mem[14][76] , \key_mem[14][75] , 
       \key_mem[14][74] , \key_mem[14][73] , \key_mem[14][72] , \key_mem[14][71] , 
       \key_mem[14][70] , \key_mem[14][69] , \key_mem[14][68] , \key_mem[14][67] , 
       \key_mem[14][66] , \key_mem[14][65] , \key_mem[14][64] , \key_mem[14][63] , 
       \key_mem[14][62] , \key_mem[14][61] , \key_mem[14][60] , \key_mem[14][59] , 
       \key_mem[14][58] , \key_mem[14][57] , \key_mem[14][56] , \key_mem[14][55] , 
       \key_mem[14][54] , \key_mem[14][53] , \key_mem[14][52] , \key_mem[14][51] , 
       \key_mem[14][50] , \key_mem[14][49] , \key_mem[14][48] , \key_mem[14][47] , 
       \key_mem[14][46] , \key_mem[14][45] , \key_mem[14][44] , \key_mem[14][43] , 
       \key_mem[14][42] , \key_mem[14][41] , \key_mem[14][40] , \key_mem[14][39] , 
       \key_mem[14][38] , \key_mem[14][37] , \key_mem[14][36] , \key_mem[14][35] , 
       \key_mem[14][34] , \key_mem[14][33] , \key_mem[14][32] , \key_mem[14][31] , 
       \key_mem[14][30] , \key_mem[14][29] , \key_mem[14][28] , \key_mem[14][27] , 
       \key_mem[14][26] , \key_mem[14][25] , \key_mem[14][24] , \key_mem[14][23] , 
       \key_mem[14][22] , \key_mem[14][21] , \key_mem[14][20] , \key_mem[14][19] , 
       \key_mem[14][18] , \key_mem[14][17] , \key_mem[14][16] , \key_mem[14][15] , 
       \key_mem[14][14] , \key_mem[14][13] , \key_mem[14][12] , \key_mem[14][11] , 
       \key_mem[14][10] , \key_mem[14][9] , \key_mem[14][8] , \key_mem[14][7] , 
       \key_mem[14][6] , \key_mem[14][5] , \key_mem[14][4] , \key_mem[14][3] , 
       \key_mem[14][2] , \key_mem[14][1] , \key_mem[14][0] , n2212, n2213, n2214, n2215, 
       n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227
       , n2228, n2229, n2230, n2242, n2243, n2276, n2277, n2278, n2282, n2283, n2284, 
       n2286, n2288, n2289, n2290, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299
       , n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
       n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322
       , n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, 
       n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345
       , n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, 
       n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368
       , n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, 
       n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391
       , n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, 
       n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414
       , n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, 
       n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437
       , n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, 
       n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460
       , n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, 
       n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483
       , n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, 
       n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506
       , n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, 
       n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529
       , n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
       n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552
       , n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, 
       n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575
       , n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, 
       n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598
       , n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, 
       n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621
       , n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, 
       n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644
       , n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, 
       n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667
       , n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, 
       n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690
       , n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, 
       n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713
       , n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
       n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736
       , n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, 
       n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759
       , n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
       n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782
       , n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, 
       n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805
       , n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, 
       n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828
       , n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
       n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851
       , n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, 
       n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874
       , n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, 
       n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897
       , n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, 
       n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920
       , n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, 
       n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943
       , n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, 
       n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966
       , n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
       n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989
       , n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
       n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012
       , n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
       n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035
       , n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, 
       n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058
       , n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, 
       n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081
       , n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, 
       n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104
       , n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, 
       n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127
       , n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, 
       n3139, n3140, n3141, n3142, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151
       , n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, 
       n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174
       , n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, 
       n3186, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198
       , n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, 
       n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221
       , n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, 
       n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244
       , n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, 
       n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267
       , n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, 
       n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291
       , n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, 
       n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314
       , n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3325, n3326, 
       n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3335, n3336, n3337, n3338, n3339
       , n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3350, n3351, 
       n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363
       , n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, 
       n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386
       , n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, 
       n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3410
       , n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, 
       n3423, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435
       , n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, 
       n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458
       , n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, 
       n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481
       , n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, 
       n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504
       , n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, 
       n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527
       , n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, 
       n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550
       , n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, 
       n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573
       , n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, 
       n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596
       , n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
       n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619
       , n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
       n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642
       , n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
       n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665
       , n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
       n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688
       , n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, 
       n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711
       , n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, 
       n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734
       , n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, 
       n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757
       , n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, 
       n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780
       , n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
       n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803
       , n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
       n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826
       , n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
       n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849
       , n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, 
       n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872
       , n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
       n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895
       , n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
       n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918
       , n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, 
       n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941
       , n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, 
       n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964
       , n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, 
       n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987
       , n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, 
       n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010
       , n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
       n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033
       , n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, 
       n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056
       , n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
       n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079
       , n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
       n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102
       , n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, 
       n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125
       , n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, 
       n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148
       , n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, 
       n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171
       , n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, 
       n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194
       , n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, 
       n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217
       , n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, 
       n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240
       , n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, 
       n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263
       , n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
       n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286
       , n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
       n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309
       , n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, 
       n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332
       , n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
       n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355
       , n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
       n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378
       , n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, 
       n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401
       , n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, 
       n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424
       , n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, 
       n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447
       , n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
       n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470
       , n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, 
       n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493
       , n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
       n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516
       , n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
       n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539
       , n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, 
       n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562
       , n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
       n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585
       , n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, 
       n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608
       , n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, 
       n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631
       , n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
       n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654
       , n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, 
       n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677
       , n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, 
       n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700
       , n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, 
       n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723
       , n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, 
       n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746
       , n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
       n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769
       , n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, 
       n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792
       , n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
       n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815
       , n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, 
       n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838
       , n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, 
       n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861
       , n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, 
       n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884
       , n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, 
       n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907
       , n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, 
       n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930
       , n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
       n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953
       , n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, 
       n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976
       , n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, 
       n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999
       , n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
       n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022
       , n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
       n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045
       , n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, 
       n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068
       , n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, 
       n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091
       , n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, 
       n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114
       , n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, 
       n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137
       , n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, 
       n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160
       , n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, 
       n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183
       , n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, 
       n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206
       , n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
       n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229
       , n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, 
       n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252
       , n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, 
       n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275
       , n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, 
       n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298
       , n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
       n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321
       , n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
       n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344
       , n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, 
       n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367
       , n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, 
       n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390
       , n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, 
       n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413
       , n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, 
       n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436
       , n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
       n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459
       , n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, 
       n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482
       , n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, 
       n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505
       , n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, 
       n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528
       , n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
       n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551
       , n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
       n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574
       , n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, 
       n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597
       , n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, 
       n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n1, n2, n3, n4, n2196, 
       n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208
       , n2209, n2210, n2211, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, 
       n2239, n2240, n2241, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252
       , n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, 
       n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275
       , n2279, n2280, n2281, n2285, n2287, n2291, n3143, n3187, n3279, n3324, n3334, 
       n3349, n3409, n3422, n3424, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624
       , n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, 
       n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647
       , n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, 
       n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670
       , n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
       n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693
       , n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
       n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716
       , n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
       n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739
       , n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, 
       n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762
       , n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, 
       n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785
       , n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, 
       n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808
       , n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, 
       n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831
       , n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
       n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854
       , n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, 
       n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877
       , n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, 
       n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900
       , n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
       n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923
       , n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, 
       n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946
       , n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
       n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969
       , n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, 
       n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992
       , n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
       n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015
       , n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, 
       n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038
       , n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
       n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061
       , n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, 
       n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084
       , n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, 
       n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107
       , n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, 
       n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130
       , n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
       n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153
       , n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, 
       n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176
       , n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
       n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199
       , n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, 
       n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222
       , n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, 
       n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245
       , n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, 
       n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268
       , n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, 
       n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291
       , n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, 
       n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314
       , n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, 
       n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337
       , n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, 
       n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360
       , n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
       n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383
       , n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, 
       n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406
       , n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
       n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429
       , n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, 
       n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452
       , n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, 
       n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475
       , n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, 
       n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498
       , n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, 
       n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521
       , n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
       n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544
       , n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, 
       n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567
       , n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, 
       n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590
       , n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
       n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613
       , n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, 
       n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636
       , n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, 
       n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659
       , n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, 
       n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682
       , n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, 
       n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705
       , n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, 
       n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728
       , n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, 
       n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751
       , n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, 
       n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774
       , n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
       n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797
       , n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, 
       n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820
       , n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
       n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843
       , n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, 
       n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866
       , n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, 
       n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889
       , n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, 
       n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912
       , n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, 
       n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935
       , n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, 
       n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958
       , n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, 
       n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981
       , n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, 
       n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004
       , n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
       n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027
       , n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, 
       n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050
       , n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
       n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073
       , n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, 
       n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096
       , n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, 
       n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119
       , n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, 
       n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142
       , n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, 
       n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165
       , n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, 
       n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188
       , n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, 
       n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211
       , n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
       n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234
       , n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, 
       n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257
       , n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, 
       n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280
       , n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
       n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303
       , n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, 
       n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326
       , n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, 
       n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349
       , n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, 
       n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372
       , n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
       n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395
       , n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, 
       n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418
       , n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, 
       n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441
       , n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, 
       n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464
       , n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, 
       n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487
       , n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, 
       n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510
       , n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, 
       n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533
       , n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, 
       n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556
       , n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, 
       n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579
       , n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, 
       n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602
       , n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
       n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7624, n7625, n7626
       , n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, 
       n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649
       , n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, 
       n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672
       , n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
       n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695
       , n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, 
       n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718
       , n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, 
       n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741
       , n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, 
       n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764
       , n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, 
       n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787
       , n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, 
       n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810
       , n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, 
       n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833
       , n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, 
       n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856
       , n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, 
       n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879
       , n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, 
       n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902
       , n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
       n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925
       , n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, 
       n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948
       , n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, 
       n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971
       , n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, 
       n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994
       , n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, 
       n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017
       , n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, 
       n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040
       , n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, 
       n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063
       , n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, 
       n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086
       , n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, 
       n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109
       , n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, 
       n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132
       , n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
       n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155
       , n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, 
       n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178
       , n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, 
       n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201
       , n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, 
       n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224
       , n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, 
       n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247
       , n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, 
       n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270
       , n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, 
       n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293
       , n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, 
       n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316
       , n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, 
       n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339
       , n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, 
       n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362
       , n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
       n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385
       , n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, 
       n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408
       , n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, 
       n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431
       , n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, 
       n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454
       , n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, 
       n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477
       , n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, 
       n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500
       , n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, 
       n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523
       , n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, 
       n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546
       , n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, 
       n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569
       , n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, 
       n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592
       , n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
       n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615
       , n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, 
       n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638
       , n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, 
       n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661
       , n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, 
       n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684
       , n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, 
       n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707
       , n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, 
       n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730
       , n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, 
       n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753
       , n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, 
       n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776
       , n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, 
       n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799
       , n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, 
       n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822
       , n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
       n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845
       , n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, 
       n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868
       , n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, 
       n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891
       , n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, 
       n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914
       , n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, 
       n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937
       , n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, 
       n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960
       , n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, 
       n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983
       , n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, 
       n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006
       , n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, 
       n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029
       , n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, 
       n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052
       , n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
       n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075
       , n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, 
       n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098
       , n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, 
       n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121
       , n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, 
       n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144
       , n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, 
       n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167
       , n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, 
       n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190
       , n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, 
       n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213
       , n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, 
       n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236
       , n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
       n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259
       , n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, 
       n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282
       , n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
       n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305
       , n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, 
       n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328
       , n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, 
       n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351
       , n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, 
       n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374
       , n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, 
       n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397
       , n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, 
       n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420
       , n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, 
       n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443
       , n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, 
       n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466
       , n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
       n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489
       , n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, 
       n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512
       , n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
       n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535
       , n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, 
       n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558
       , n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, 
       n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581
       , n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, 
       n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604
       , n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, 
       n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627
       , n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, 
       n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650
       , n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, 
       n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673
       , n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, 
       n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696
       , n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, 
       n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719
       , n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, 
       n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742
       , n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
       n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765
       , n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
       n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, clk_buf_net0, 
       clk_buf_net1, clk_buf_net2, clk_buf_net3, clk_buf_net4, clk_buf_net5, clk_buf_net6
       , clk_buf_net7, test_se_buf_net0, test_se_buf_net1, test_se_buf_net2, 
       test_se_buf_net3, test_se_buf_net4, test_se_buf_net5, test_se_buf_net6, 
       test_se_buf_net7;
wire [7:0] rcon_reg;
wire [127:0] prev_key0_reg;
wire [127:32] prev_key1_reg;
wire [2:0] key_mem_ctrl_reg;
wire [3:0] round_ctr_reg;
   assign N28 = round[0];
   assign N29 = round[1];
   assign N30 = round[2];
   assign N31 = round[3];
   assign test_so1 = \key_mem[4][77] ;
   assign test_so2 = \key_mem[12][49] ;
   assign test_so3 = n2212;
   SDFFARX1 \key_mem_ctrl_reg_reg[0]  (.D(n5616), .SI(test_si1), .SE(test_se), .CLK(clk), .
          RSTB(n7495), .Q(key_mem_ctrl_reg[0]), .QN(n2243));
   SDFFARX1 \round_ctr_reg_reg[1]  (.D(n5613), .SI(round_ctr_reg[0]), .SE(test_se), .CLK(
          clk), .RSTB(n7495), .Q(round_ctr_reg[1]), .QN(n2213));
   SDFFARX1 \round_ctr_reg_reg[3]  (.D(n5611), .SI(n7624), .SE(test_se), .CLK(clk), .RSTB(
          n7495), .Q(round_ctr_reg[3]), .QN(n2212));
   SDFFARX1 \rcon_reg_reg[0]  (.D(n5609), .SI(n7634), .SE(test_se), .CLK(clk), .RSTB(n7495)
          , .Q(rcon_reg[0]), .QN(n7633));
   SDFFARX1 \rcon_reg_reg[1]  (.D(n5610), .SI(n7633), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[1]), .QN(n7632));
   SDFFARX1 \rcon_reg_reg[2]  (.D(n5608), .SI(n7632), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[2]), .QN(n7631));
   SDFFARX1 \rcon_reg_reg[3]  (.D(n5607), .SI(n7631), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[3]), .QN(n7630));
   SDFFARX1 \rcon_reg_reg[4]  (.D(n5606), .SI(n7630), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[4]), .QN(n7629));
   SDFFARX1 \rcon_reg_reg[5]  (.D(n5605), .SI(n7629), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[5]), .QN(n7628));
   SDFFARX1 \rcon_reg_reg[6]  (.D(n5604), .SI(n7628), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[6]), .QN(n7627));
   SDFFARX1 \rcon_reg_reg[7]  (.D(n5603), .SI(n7627), .SE(test_se), .CLK(clk), .RSTB(n7494)
          , .Q(rcon_reg[7]), .QN(n7626));
   SDFFARX1 ready_reg_reg (.D(n5602), .SI(n7626), .SE(test_se), .CLK(clk), .RSTB(n7494), .
          Q(ready), .QN(n7625));
   SDFFARX1 \prev_key1_reg_reg[127]  (.D(n5346), .SI(n7635), .SE(test_se), .CLK(clk), .
          RSTB(n7494), .Q(prev_key1_reg[127]), .QN(n7634));
   SDFFARX1 \prev_key0_reg_reg[127]  (.D(n5473), .SI(prev_key0_reg[126]), .SE(test_se), .
          CLK(clk), .RSTB(n7494), .Q(prev_key0_reg[127]), .QN(n2215));
   SDFFARX1 \key_mem_reg[0][127]  (.D(n3426), .SI(n9659), .SE(test_se), .CLK(clk), .RSTB(
          n7494), .Q(\key_mem[0][127] ), .QN(n9658));
   SDFFARX1 \key_mem_reg[1][127]  (.D(n3427), .SI(n9531), .SE(test_se), .CLK(clk), .RSTB(
          n7494), .Q(\key_mem[1][127] ), .QN(n9530));
   SDFFARX1 \key_mem_reg[2][127]  (.D(n3428), .SI(n9403), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[2][127] ), .QN(n9402));
   SDFFARX1 \key_mem_reg[3][127]  (.D(n3429), .SI(n9275), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[3][127] ), .QN(n9274));
   SDFFARX1 \key_mem_reg[4][127]  (.D(n3430), .SI(n9148), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[4][127] ), .QN(n9147));
   SDFFARX1 \key_mem_reg[5][127]  (.D(n3431), .SI(n9020), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[5][127] ), .QN(n9019));
   SDFFARX1 \key_mem_reg[6][127]  (.D(n3432), .SI(n8892), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[6][127] ), .QN(n8891));
   SDFFARX1 \key_mem_reg[7][127]  (.D(n3433), .SI(n8764), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[7][127] ), .QN(n8763));
   SDFFARX1 \key_mem_reg[8][127]  (.D(n3434), .SI(n8636), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[8][127] ), .QN(n8635));
   SDFFARX1 \key_mem_reg[9][127]  (.D(n3435), .SI(n8508), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[9][127] ), .QN(n8507));
   SDFFARX1 \key_mem_reg[10][127]  (.D(n3436), .SI(n8380), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[10][127] ), .QN(n8379));
   SDFFARX1 \key_mem_reg[11][127]  (.D(n3437), .SI(n8252), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[11][127] ), .QN(n8251));
   SDFFARX1 \key_mem_reg[12][127]  (.D(n3438), .SI(n8125), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[12][127] ), .QN(n8124));
   SDFFARX1 \key_mem_reg[13][127]  (.D(n3439), .SI(n7997), .SE(test_se), .CLK(clk), .RSTB(
          n7493), .Q(\key_mem[13][127] ), .QN(n7996));
   SDFFARX1 \key_mem_reg[14][127]  (.D(n3440), .SI(n7869), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[14][127] ), .QN(n7868));
   SDFFARX1 \prev_key1_reg_reg[126]  (.D(n5347), .SI(n7636), .SE(test_se), .CLK(clk), .
          RSTB(n7492), .Q(prev_key1_reg[126]), .QN(n7635));
   SDFFARX1 \prev_key0_reg_reg[126]  (.D(n5474), .SI(prev_key0_reg[125]), .SE(test_se), .
          CLK(clk), .RSTB(n7492), .Q(prev_key0_reg[126]), .QN(n2216));
   SDFFARX1 \key_mem_reg[0][126]  (.D(n3441), .SI(n9660), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[0][126] ), .QN(n9659));
   SDFFARX1 \key_mem_reg[1][126]  (.D(n3442), .SI(n9532), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[1][126] ), .QN(n9531));
   SDFFARX1 \key_mem_reg[2][126]  (.D(n3443), .SI(n9404), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[2][126] ), .QN(n9403));
   SDFFARX1 \key_mem_reg[3][126]  (.D(n3444), .SI(n9276), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[3][126] ), .QN(n9275));
   SDFFARX1 \key_mem_reg[4][126]  (.D(n3445), .SI(n9149), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[4][126] ), .QN(n9148));
   SDFFARX1 \key_mem_reg[5][126]  (.D(n3446), .SI(n9021), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[5][126] ), .QN(n9020));
   SDFFARX1 \key_mem_reg[6][126]  (.D(n3447), .SI(n8893), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[6][126] ), .QN(n8892));
   SDFFARX1 \key_mem_reg[7][126]  (.D(n3448), .SI(n8765), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[7][126] ), .QN(n8764));
   SDFFARX1 \key_mem_reg[8][126]  (.D(n3449), .SI(n8637), .SE(test_se), .CLK(clk), .RSTB(
          n7492), .Q(\key_mem[8][126] ), .QN(n8636));
   SDFFARX1 \key_mem_reg[9][126]  (.D(n3450), .SI(n8509), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[9][126] ), .QN(n8508));
   SDFFARX1 \key_mem_reg[10][126]  (.D(n3451), .SI(n8381), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[10][126] ), .QN(n8380));
   SDFFARX1 \key_mem_reg[11][126]  (.D(n3452), .SI(n8253), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[11][126] ), .QN(n8252));
   SDFFARX1 \key_mem_reg[12][126]  (.D(n3453), .SI(n8126), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[12][126] ), .QN(n8125));
   SDFFARX1 \key_mem_reg[13][126]  (.D(n3454), .SI(n7998), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[13][126] ), .QN(n7997));
   SDFFARX1 \key_mem_reg[14][126]  (.D(n3455), .SI(n7870), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[14][126] ), .QN(n7869));
   SDFFARX1 \prev_key1_reg_reg[125]  (.D(n5348), .SI(n7637), .SE(test_se), .CLK(clk), .
          RSTB(n7491), .Q(prev_key1_reg[125]), .QN(n7636));
   SDFFARX1 \prev_key0_reg_reg[125]  (.D(n5475), .SI(prev_key0_reg[124]), .SE(test_se), .
          CLK(clk), .RSTB(n7491), .Q(prev_key0_reg[125]), .QN(n2217));
   SDFFARX1 \key_mem_reg[0][125]  (.D(n3456), .SI(n9661), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[0][125] ), .QN(n9660));
   SDFFARX1 \key_mem_reg[1][125]  (.D(n3457), .SI(n9533), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[1][125] ), .QN(n9532));
   SDFFARX1 \key_mem_reg[2][125]  (.D(n3458), .SI(n9405), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[2][125] ), .QN(n9404));
   SDFFARX1 \key_mem_reg[3][125]  (.D(n3459), .SI(n9277), .SE(test_se), .CLK(clk), .RSTB(
          n7491), .Q(\key_mem[3][125] ), .QN(n9276));
   SDFFARX1 \key_mem_reg[4][125]  (.D(n3460), .SI(n9150), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[4][125] ), .QN(n9149));
   SDFFARX1 \key_mem_reg[5][125]  (.D(n3461), .SI(n9022), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[5][125] ), .QN(n9021));
   SDFFARX1 \key_mem_reg[6][125]  (.D(n3462), .SI(n8894), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[6][125] ), .QN(n8893));
   SDFFARX1 \key_mem_reg[7][125]  (.D(n3463), .SI(n8766), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[7][125] ), .QN(n8765));
   SDFFARX1 \key_mem_reg[8][125]  (.D(n3464), .SI(n8638), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[8][125] ), .QN(n8637));
   SDFFARX1 \key_mem_reg[9][125]  (.D(n3465), .SI(n8510), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[9][125] ), .QN(n8509));
   SDFFARX1 \key_mem_reg[10][125]  (.D(n3466), .SI(n8382), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[10][125] ), .QN(n8381));
   SDFFARX1 \key_mem_reg[11][125]  (.D(n3467), .SI(n8254), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[11][125] ), .QN(n8253));
   SDFFARX1 \key_mem_reg[12][125]  (.D(n3468), .SI(n8127), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[12][125] ), .QN(n8126));
   SDFFARX1 \key_mem_reg[13][125]  (.D(n3469), .SI(n7999), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[13][125] ), .QN(n7998));
   SDFFARX1 \key_mem_reg[14][125]  (.D(n3470), .SI(n7871), .SE(test_se), .CLK(clk), .RSTB(
          n7490), .Q(\key_mem[14][125] ), .QN(n7870));
   SDFFARX1 \prev_key1_reg_reg[124]  (.D(n5349), .SI(n7638), .SE(test_se), .CLK(clk), .
          RSTB(n7490), .Q(prev_key1_reg[124]), .QN(n7637));
   SDFFARX1 \prev_key0_reg_reg[124]  (.D(n5476), .SI(prev_key0_reg[123]), .SE(test_se), .
          CLK(clk), .RSTB(n7489), .Q(prev_key0_reg[124]), .QN(n2218));
   SDFFARX1 \key_mem_reg[0][124]  (.D(n3471), .SI(n9662), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[0][124] ), .QN(n9661));
   SDFFARX1 \key_mem_reg[1][124]  (.D(n3472), .SI(n9534), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[1][124] ), .QN(n9533));
   SDFFARX1 \key_mem_reg[2][124]  (.D(n3473), .SI(n9406), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[2][124] ), .QN(n9405));
   SDFFARX1 \key_mem_reg[3][124]  (.D(n3474), .SI(n9278), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[3][124] ), .QN(n9277));
   SDFFARX1 \key_mem_reg[4][124]  (.D(n3475), .SI(n9151), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[4][124] ), .QN(n9150));
   SDFFARX1 \key_mem_reg[5][124]  (.D(n3476), .SI(n9023), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[5][124] ), .QN(n9022));
   SDFFARX1 \key_mem_reg[6][124]  (.D(n3477), .SI(n8895), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[6][124] ), .QN(n8894));
   SDFFARX1 \key_mem_reg[7][124]  (.D(n3478), .SI(n8767), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[7][124] ), .QN(n8766));
   SDFFARX1 \key_mem_reg[8][124]  (.D(n3479), .SI(n8639), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[8][124] ), .QN(n8638));
   SDFFARX1 \key_mem_reg[9][124]  (.D(n3480), .SI(n8511), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[9][124] ), .QN(n8510));
   SDFFARX1 \key_mem_reg[10][124]  (.D(n3481), .SI(n8383), .SE(test_se), .CLK(clk), .RSTB(
          n7489), .Q(\key_mem[10][124] ), .QN(n8382));
   SDFFARX1 \key_mem_reg[11][124]  (.D(n3482), .SI(n8255), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[11][124] ), .QN(n8254));
   SDFFARX1 \key_mem_reg[12][124]  (.D(n3483), .SI(n8128), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[12][124] ), .QN(n8127));
   SDFFARX1 \key_mem_reg[13][124]  (.D(n3484), .SI(n8000), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[13][124] ), .QN(n7999));
   SDFFARX1 \key_mem_reg[14][124]  (.D(n3485), .SI(n7872), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[14][124] ), .QN(n7871));
   SDFFARX1 \prev_key1_reg_reg[123]  (.D(n5350), .SI(n7639), .SE(test_se), .CLK(clk), .
          RSTB(n7488), .Q(prev_key1_reg[123]), .QN(n7638));
   SDFFARX1 \prev_key0_reg_reg[123]  (.D(n5477), .SI(prev_key0_reg[122]), .SE(test_se), .
          CLK(clk), .RSTB(n7488), .Q(prev_key0_reg[123]), .QN(n2219));
   SDFFARX1 \key_mem_reg[0][123]  (.D(n3486), .SI(n9663), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[0][123] ), .QN(n9662));
   SDFFARX1 \key_mem_reg[1][123]  (.D(n3487), .SI(n9535), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[1][123] ), .QN(n9534));
   SDFFARX1 \key_mem_reg[2][123]  (.D(n3488), .SI(n9407), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[2][123] ), .QN(n9406));
   SDFFARX1 \key_mem_reg[3][123]  (.D(n3489), .SI(n9279), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[3][123] ), .QN(n9278));
   SDFFARX1 \key_mem_reg[4][123]  (.D(n3490), .SI(n9152), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[4][123] ), .QN(n9151));
   SDFFARX1 \key_mem_reg[5][123]  (.D(n3491), .SI(n9024), .SE(test_se), .CLK(clk), .RSTB(
          n7488), .Q(\key_mem[5][123] ), .QN(n9023));
   SDFFARX1 \key_mem_reg[6][123]  (.D(n3492), .SI(n8896), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[6][123] ), .QN(n8895));
   SDFFARX1 \key_mem_reg[7][123]  (.D(n3493), .SI(n8768), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[7][123] ), .QN(n8767));
   SDFFARX1 \key_mem_reg[8][123]  (.D(n3494), .SI(n8640), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[8][123] ), .QN(n8639));
   SDFFARX1 \key_mem_reg[9][123]  (.D(n3495), .SI(n8512), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[9][123] ), .QN(n8511));
   SDFFARX1 \key_mem_reg[10][123]  (.D(n3496), .SI(n8384), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[10][123] ), .QN(n8383));
   SDFFARX1 \key_mem_reg[11][123]  (.D(n3497), .SI(n8256), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[11][123] ), .QN(n8255));
   SDFFARX1 \key_mem_reg[12][123]  (.D(n3498), .SI(n8129), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[12][123] ), .QN(n8128));
   SDFFARX1 \key_mem_reg[13][123]  (.D(n3499), .SI(n8001), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[13][123] ), .QN(n8000));
   SDFFARX1 \key_mem_reg[14][123]  (.D(n3500), .SI(n7873), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[14][123] ), .QN(n7872));
   SDFFARX1 \prev_key1_reg_reg[122]  (.D(n5351), .SI(n7640), .SE(test_se), .CLK(clk), .
          RSTB(n7487), .Q(prev_key1_reg[122]), .QN(n7639));
   SDFFARX1 \prev_key0_reg_reg[122]  (.D(n5478), .SI(prev_key0_reg[121]), .SE(test_se), .
          CLK(clk), .RSTB(n7487), .Q(prev_key0_reg[122]), .QN(n2220));
   SDFFARX1 \key_mem_reg[0][122]  (.D(n3501), .SI(n9664), .SE(test_se), .CLK(clk), .RSTB(
          n7487), .Q(\key_mem[0][122] ), .QN(n9663));
   SDFFARX1 \key_mem_reg[1][122]  (.D(n3502), .SI(n9536), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[1][122] ), .QN(n9535));
   SDFFARX1 \key_mem_reg[2][122]  (.D(n3503), .SI(n9408), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[2][122] ), .QN(n9407));
   SDFFARX1 \key_mem_reg[3][122]  (.D(n3504), .SI(n9280), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[3][122] ), .QN(n9279));
   SDFFARX1 \key_mem_reg[4][122]  (.D(n3505), .SI(n9153), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[4][122] ), .QN(n9152));
   SDFFARX1 \key_mem_reg[5][122]  (.D(n3506), .SI(n9025), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[5][122] ), .QN(n9024));
   SDFFARX1 \key_mem_reg[6][122]  (.D(n3507), .SI(n8897), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[6][122] ), .QN(n8896));
   SDFFARX1 \key_mem_reg[7][122]  (.D(n3508), .SI(n8769), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[7][122] ), .QN(n8768));
   SDFFARX1 \key_mem_reg[8][122]  (.D(n3509), .SI(n8641), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[8][122] ), .QN(n8640));
   SDFFARX1 \key_mem_reg[9][122]  (.D(n3510), .SI(n8513), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[9][122] ), .QN(n8512));
   SDFFARX1 \key_mem_reg[10][122]  (.D(n3511), .SI(n8385), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[10][122] ), .QN(n8384));
   SDFFARX1 \key_mem_reg[11][122]  (.D(n3512), .SI(n8257), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[11][122] ), .QN(n8256));
   SDFFARX1 \key_mem_reg[12][122]  (.D(n3513), .SI(n8130), .SE(test_se), .CLK(clk), .RSTB(
          n7486), .Q(\key_mem[12][122] ), .QN(n8129));
   SDFFARX1 \key_mem_reg[13][122]  (.D(n3514), .SI(n8002), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[13][122] ), .QN(n8001));
   SDFFARX1 \key_mem_reg[14][122]  (.D(n3515), .SI(n7874), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[14][122] ), .QN(n7873));
   SDFFARX1 \prev_key1_reg_reg[121]  (.D(n5352), .SI(n4), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(prev_key1_reg[121]), .QN(n7640));
   SDFFARX1 \prev_key0_reg_reg[121]  (.D(n5479), .SI(prev_key0_reg[120]), .SE(test_se), .
          CLK(clk), .RSTB(n7485), .Q(prev_key0_reg[121]), .QN(n2221));
   SDFFARX1 \key_mem_reg[0][121]  (.D(n3516), .SI(n9665), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[0][121] ), .QN(n9664));
   SDFFARX1 \key_mem_reg[1][121]  (.D(n3517), .SI(n9537), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[1][121] ), .QN(n9536));
   SDFFARX1 \key_mem_reg[2][121]  (.D(n3518), .SI(n9409), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[2][121] ), .QN(n9408));
   SDFFARX1 \key_mem_reg[3][121]  (.D(n3519), .SI(n9281), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[3][121] ), .QN(n9280));
   SDFFARX1 \key_mem_reg[4][121]  (.D(n3520), .SI(n9154), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[4][121] ), .QN(n9153));
   SDFFARX1 \key_mem_reg[5][121]  (.D(n3521), .SI(n9026), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[5][121] ), .QN(n9025));
   SDFFARX1 \key_mem_reg[6][121]  (.D(n3522), .SI(n8898), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[6][121] ), .QN(n8897));
   SDFFARX1 \key_mem_reg[7][121]  (.D(n3523), .SI(n8770), .SE(test_se), .CLK(clk), .RSTB(
          n7485), .Q(\key_mem[7][121] ), .QN(n8769));
   SDFFARX1 \key_mem_reg[8][121]  (.D(n3524), .SI(n8642), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[8][121] ), .QN(n8641));
   SDFFARX1 \key_mem_reg[9][121]  (.D(n3525), .SI(n8514), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[9][121] ), .QN(n8513));
   SDFFARX1 \key_mem_reg[10][121]  (.D(n3526), .SI(n8386), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[10][121] ), .QN(n8385));
   SDFFARX1 \key_mem_reg[11][121]  (.D(n3527), .SI(n8258), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[11][121] ), .QN(n8257));
   SDFFARX1 \key_mem_reg[12][121]  (.D(n3528), .SI(n8131), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[12][121] ), .QN(n8130));
   SDFFARX1 \key_mem_reg[13][121]  (.D(n3529), .SI(n8003), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[13][121] ), .QN(n8002));
   SDFFARX1 \key_mem_reg[14][121]  (.D(n3530), .SI(n7875), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[14][121] ), .QN(n7874));
   SDFFARX1 \prev_key1_reg_reg[120]  (.D(n5353), .SI(n7641), .SE(test_se), .CLK(clk), .
          RSTB(n7484), .Q(prev_key1_reg[120]), .QN(n4));
   SDFFARX1 \prev_key0_reg_reg[120]  (.D(n5480), .SI(prev_key0_reg[119]), .SE(test_se), .
          CLK(clk), .RSTB(n7484), .Q(prev_key0_reg[120]), .QN(n2222));
   SDFFARX1 \key_mem_reg[0][120]  (.D(n3531), .SI(n9666), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[0][120] ), .QN(n9665));
   SDFFARX1 \key_mem_reg[1][120]  (.D(n3532), .SI(n9538), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[1][120] ), .QN(n9537));
   SDFFARX1 \key_mem_reg[2][120]  (.D(n3533), .SI(n9410), .SE(test_se), .CLK(clk), .RSTB(
          n7484), .Q(\key_mem[2][120] ), .QN(n9409));
   SDFFARX1 \key_mem_reg[3][120]  (.D(n3534), .SI(n9282), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[3][120] ), .QN(n9281));
   SDFFARX1 \key_mem_reg[4][120]  (.D(n3535), .SI(n9155), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[4][120] ), .QN(n9154));
   SDFFARX1 \key_mem_reg[5][120]  (.D(n3536), .SI(n9027), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[5][120] ), .QN(n9026));
   SDFFARX1 \key_mem_reg[6][120]  (.D(n3537), .SI(n8899), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[6][120] ), .QN(n8898));
   SDFFARX1 \key_mem_reg[7][120]  (.D(n3538), .SI(n8771), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[7][120] ), .QN(n8770));
   SDFFARX1 \key_mem_reg[8][120]  (.D(n3539), .SI(n8643), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[8][120] ), .QN(n8642));
   SDFFARX1 \key_mem_reg[9][120]  (.D(n3540), .SI(n8515), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[9][120] ), .QN(n8514));
   SDFFARX1 \key_mem_reg[10][120]  (.D(n3541), .SI(n8387), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[10][120] ), .QN(n8386));
   SDFFARX1 \key_mem_reg[11][120]  (.D(n3542), .SI(n8259), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[11][120] ), .QN(n8258));
   SDFFARX1 \key_mem_reg[12][120]  (.D(n3543), .SI(n8132), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[12][120] ), .QN(n8131));
   SDFFARX1 \key_mem_reg[13][120]  (.D(n3544), .SI(n8004), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[13][120] ), .QN(n8003));
   SDFFARX1 \key_mem_reg[14][120]  (.D(n3545), .SI(n7876), .SE(test_se), .CLK(clk), .RSTB(
          n7483), .Q(\key_mem[14][120] ), .QN(n7875));
   SDFFARX1 \prev_key1_reg_reg[119]  (.D(n5354), .SI(n7642), .SE(test_se), .CLK(clk), .
          RSTB(n7482), .Q(prev_key1_reg[119]), .QN(n7641));
   SDFFARX1 \prev_key0_reg_reg[119]  (.D(n5481), .SI(prev_key0_reg[118]), .SE(test_se), .
          CLK(clk), .RSTB(n7482), .Q(prev_key0_reg[119]), .QN(n2223));
   SDFFARX1 \key_mem_reg[0][119]  (.D(n3546), .SI(n9667), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[0][119] ), .QN(n9666));
   SDFFARX1 \key_mem_reg[1][119]  (.D(n3547), .SI(n9539), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[1][119] ), .QN(n9538));
   SDFFARX1 \key_mem_reg[2][119]  (.D(n3548), .SI(n9411), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[2][119] ), .QN(n9410));
   SDFFARX1 \key_mem_reg[3][119]  (.D(n3549), .SI(n9283), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[3][119] ), .QN(n9282));
   SDFFARX1 \key_mem_reg[4][119]  (.D(n3550), .SI(n9156), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[4][119] ), .QN(n9155));
   SDFFARX1 \key_mem_reg[5][119]  (.D(n3551), .SI(n9028), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[5][119] ), .QN(n9027));
   SDFFARX1 \key_mem_reg[6][119]  (.D(n3552), .SI(n8900), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[6][119] ), .QN(n8899));
   SDFFARX1 \key_mem_reg[7][119]  (.D(n3553), .SI(n8772), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[7][119] ), .QN(n8771));
   SDFFARX1 \key_mem_reg[8][119]  (.D(n3554), .SI(n8644), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[8][119] ), .QN(n8643));
   SDFFARX1 \key_mem_reg[9][119]  (.D(n3555), .SI(n8516), .SE(test_se), .CLK(clk), .RSTB(
          n7482), .Q(\key_mem[9][119] ), .QN(n8515));
   SDFFARX1 \key_mem_reg[10][119]  (.D(n3556), .SI(n8388), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[10][119] ), .QN(n8387));
   SDFFARX1 \key_mem_reg[11][119]  (.D(n3557), .SI(n8260), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[11][119] ), .QN(n8259));
   SDFFARX1 \key_mem_reg[12][119]  (.D(n3558), .SI(n8133), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[12][119] ), .QN(n8132));
   SDFFARX1 \key_mem_reg[13][119]  (.D(n3559), .SI(n8005), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[13][119] ), .QN(n8004));
   SDFFARX1 \key_mem_reg[14][119]  (.D(n3560), .SI(n7877), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[14][119] ), .QN(n7876));
   SDFFARX1 \prev_key1_reg_reg[118]  (.D(n5355), .SI(n7643), .SE(test_se), .CLK(clk), .
          RSTB(n7481), .Q(prev_key1_reg[118]), .QN(n7642));
   SDFFARX1 \prev_key0_reg_reg[118]  (.D(n5482), .SI(prev_key0_reg[117]), .SE(test_se), .
          CLK(clk), .RSTB(n7481), .Q(prev_key0_reg[118]), .QN(n2224));
   SDFFARX1 \key_mem_reg[0][118]  (.D(n3561), .SI(n9668), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[0][118] ), .QN(n9667));
   SDFFARX1 \key_mem_reg[1][118]  (.D(n3562), .SI(n9540), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[1][118] ), .QN(n9539));
   SDFFARX1 \key_mem_reg[2][118]  (.D(n3563), .SI(n9412), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[2][118] ), .QN(n9411));
   SDFFARX1 \key_mem_reg[3][118]  (.D(n3564), .SI(n9284), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[3][118] ), .QN(n9283));
   SDFFARX1 \key_mem_reg[4][118]  (.D(n3565), .SI(n9157), .SE(test_se), .CLK(clk), .RSTB(
          n7481), .Q(\key_mem[4][118] ), .QN(n9156));
   SDFFARX1 \key_mem_reg[5][118]  (.D(n3566), .SI(n9029), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[5][118] ), .QN(n9028));
   SDFFARX1 \key_mem_reg[6][118]  (.D(n3567), .SI(n8901), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[6][118] ), .QN(n8900));
   SDFFARX1 \key_mem_reg[7][118]  (.D(n3568), .SI(n8773), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[7][118] ), .QN(n8772));
   SDFFARX1 \key_mem_reg[8][118]  (.D(n3569), .SI(n8645), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[8][118] ), .QN(n8644));
   SDFFARX1 \key_mem_reg[9][118]  (.D(n3570), .SI(n8517), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[9][118] ), .QN(n8516));
   SDFFARX1 \key_mem_reg[10][118]  (.D(n3571), .SI(n8389), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[10][118] ), .QN(n8388));
   SDFFARX1 \key_mem_reg[11][118]  (.D(n3572), .SI(n8261), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[11][118] ), .QN(n8260));
   SDFFARX1 \key_mem_reg[12][118]  (.D(n3573), .SI(n8134), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[12][118] ), .QN(n8133));
   SDFFARX1 \key_mem_reg[13][118]  (.D(n3574), .SI(n8006), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[13][118] ), .QN(n8005));
   SDFFARX1 \key_mem_reg[14][118]  (.D(n3575), .SI(n7878), .SE(test_se), .CLK(clk), .RSTB(
          n7480), .Q(\key_mem[14][118] ), .QN(n7877));
   SDFFARX1 \prev_key1_reg_reg[117]  (.D(n5356), .SI(n7644), .SE(test_se), .CLK(clk), .
          RSTB(n7480), .Q(prev_key1_reg[117]), .QN(n7643));
   SDFFARX1 \prev_key0_reg_reg[117]  (.D(n5483), .SI(prev_key0_reg[116]), .SE(test_se), .
          CLK(clk), .RSTB(n7480), .Q(prev_key0_reg[117]), .QN(n2225));
   SDFFARX1 \key_mem_reg[0][117]  (.D(n3576), .SI(n9669), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[0][117] ), .QN(n9668));
   SDFFARX1 \key_mem_reg[1][117]  (.D(n3577), .SI(n9541), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[1][117] ), .QN(n9540));
   SDFFARX1 \key_mem_reg[2][117]  (.D(n3578), .SI(n9413), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[2][117] ), .QN(n9412));
   SDFFARX1 \key_mem_reg[3][117]  (.D(n3579), .SI(n9285), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[3][117] ), .QN(n9284));
   SDFFARX1 \key_mem_reg[4][117]  (.D(n3580), .SI(n9158), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[4][117] ), .QN(n9157));
   SDFFARX1 \key_mem_reg[5][117]  (.D(n3581), .SI(n9030), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[5][117] ), .QN(n9029));
   SDFFARX1 \key_mem_reg[6][117]  (.D(n3582), .SI(n8902), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[6][117] ), .QN(n8901));
   SDFFARX1 \key_mem_reg[7][117]  (.D(n3583), .SI(n8774), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[7][117] ), .QN(n8773));
   SDFFARX1 \key_mem_reg[8][117]  (.D(n3584), .SI(n8646), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[8][117] ), .QN(n8645));
   SDFFARX1 \key_mem_reg[9][117]  (.D(n3585), .SI(n8518), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[9][117] ), .QN(n8517));
   SDFFARX1 \key_mem_reg[10][117]  (.D(n3586), .SI(n8390), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[10][117] ), .QN(n8389));
   SDFFARX1 \key_mem_reg[11][117]  (.D(n3587), .SI(n8262), .SE(test_se), .CLK(clk), .RSTB(
          n7479), .Q(\key_mem[11][117] ), .QN(n8261));
   SDFFARX1 \key_mem_reg[12][117]  (.D(n3588), .SI(n8135), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[12][117] ), .QN(n8134));
   SDFFARX1 \key_mem_reg[13][117]  (.D(n3589), .SI(n8007), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[13][117] ), .QN(n8006));
   SDFFARX1 \key_mem_reg[14][117]  (.D(n3590), .SI(n7879), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[14][117] ), .QN(n7878));
   SDFFARX1 \prev_key1_reg_reg[116]  (.D(n5357), .SI(n7645), .SE(test_se), .CLK(clk), .
          RSTB(n7478), .Q(prev_key1_reg[116]), .QN(n7644));
   SDFFARX1 \prev_key0_reg_reg[116]  (.D(n5484), .SI(prev_key0_reg[115]), .SE(test_se), .
          CLK(clk), .RSTB(n7478), .Q(prev_key0_reg[116]), .QN(n2226));
   SDFFARX1 \key_mem_reg[0][116]  (.D(n3591), .SI(n9670), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[0][116] ), .QN(n9669));
   SDFFARX1 \key_mem_reg[1][116]  (.D(n3592), .SI(n9542), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[1][116] ), .QN(n9541));
   SDFFARX1 \key_mem_reg[2][116]  (.D(n3593), .SI(n9414), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[2][116] ), .QN(n9413));
   SDFFARX1 \key_mem_reg[3][116]  (.D(n3594), .SI(n9286), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[3][116] ), .QN(n9285));
   SDFFARX1 \key_mem_reg[4][116]  (.D(n3595), .SI(n9159), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[4][116] ), .QN(n9158));
   SDFFARX1 \key_mem_reg[5][116]  (.D(n3596), .SI(n9031), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[5][116] ), .QN(n9030));
   SDFFARX1 \key_mem_reg[6][116]  (.D(n3597), .SI(n8903), .SE(test_se), .CLK(clk), .RSTB(
          n7478), .Q(\key_mem[6][116] ), .QN(n8902));
   SDFFARX1 \key_mem_reg[7][116]  (.D(n3598), .SI(n8775), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[7][116] ), .QN(n8774));
   SDFFARX1 \key_mem_reg[8][116]  (.D(n3599), .SI(n8647), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[8][116] ), .QN(n8646));
   SDFFARX1 \key_mem_reg[9][116]  (.D(n3600), .SI(n8519), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[9][116] ), .QN(n8518));
   SDFFARX1 \key_mem_reg[10][116]  (.D(n3601), .SI(n8391), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[10][116] ), .QN(n8390));
   SDFFARX1 \key_mem_reg[11][116]  (.D(n3602), .SI(n8263), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[11][116] ), .QN(n8262));
   SDFFARX1 \key_mem_reg[12][116]  (.D(n3603), .SI(n8136), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[12][116] ), .QN(n8135));
   SDFFARX1 \key_mem_reg[13][116]  (.D(n3604), .SI(n8008), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[13][116] ), .QN(n8007));
   SDFFARX1 \key_mem_reg[14][116]  (.D(n3605), .SI(n7880), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[14][116] ), .QN(n7879));
   SDFFARX1 \prev_key1_reg_reg[115]  (.D(n5358), .SI(n7646), .SE(test_se), .CLK(clk), .
          RSTB(n7477), .Q(prev_key1_reg[115]), .QN(n7645));
   SDFFARX1 \prev_key0_reg_reg[115]  (.D(n5485), .SI(prev_key0_reg[114]), .SE(test_se), .
          CLK(clk), .RSTB(n7477), .Q(prev_key0_reg[115]), .QN(n2227));
   SDFFARX1 \key_mem_reg[0][115]  (.D(n3606), .SI(n9671), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[0][115] ), .QN(n9670));
   SDFFARX1 \key_mem_reg[1][115]  (.D(n3607), .SI(n9543), .SE(test_se), .CLK(clk), .RSTB(
          n7477), .Q(\key_mem[1][115] ), .QN(n9542));
   SDFFARX1 \key_mem_reg[2][115]  (.D(n3608), .SI(n9415), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[2][115] ), .QN(n9414));
   SDFFARX1 \key_mem_reg[3][115]  (.D(n3609), .SI(n9287), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[3][115] ), .QN(n9286));
   SDFFARX1 \key_mem_reg[4][115]  (.D(n3610), .SI(n9160), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[4][115] ), .QN(n9159));
   SDFFARX1 \key_mem_reg[5][115]  (.D(n3611), .SI(n9032), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[5][115] ), .QN(n9031));
   SDFFARX1 \key_mem_reg[6][115]  (.D(n3612), .SI(n8904), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[6][115] ), .QN(n8903));
   SDFFARX1 \key_mem_reg[7][115]  (.D(n3613), .SI(n8776), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[7][115] ), .QN(n8775));
   SDFFARX1 \key_mem_reg[8][115]  (.D(n3614), .SI(n8648), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[8][115] ), .QN(n8647));
   SDFFARX1 \key_mem_reg[9][115]  (.D(n3615), .SI(n8520), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[9][115] ), .QN(n8519));
   SDFFARX1 \key_mem_reg[10][115]  (.D(n3616), .SI(n8392), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[10][115] ), .QN(n8391));
   SDFFARX1 \key_mem_reg[11][115]  (.D(n3617), .SI(n8264), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[11][115] ), .QN(n8263));
   SDFFARX1 \key_mem_reg[12][115]  (.D(n3618), .SI(n8137), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[12][115] ), .QN(n8136));
   SDFFARX1 \key_mem_reg[13][115]  (.D(n3619), .SI(n8009), .SE(test_se), .CLK(clk), .RSTB(
          n7476), .Q(\key_mem[13][115] ), .QN(n8008));
   SDFFARX1 \key_mem_reg[14][115]  (.D(n3620), .SI(n7881), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[14][115] ), .QN(n7880));
   SDFFARX1 \prev_key1_reg_reg[114]  (.D(n5359), .SI(n7647), .SE(test_se), .CLK(clk), .
          RSTB(n7475), .Q(prev_key1_reg[114]), .QN(n7646));
   SDFFARX1 \prev_key0_reg_reg[114]  (.D(n5486), .SI(prev_key0_reg[113]), .SE(test_se), .
          CLK(clk), .RSTB(n7475), .Q(prev_key0_reg[114]), .QN(n2228));
   SDFFARX1 \key_mem_reg[0][114]  (.D(n3621), .SI(n9672), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[0][114] ), .QN(n9671));
   SDFFARX1 \key_mem_reg[1][114]  (.D(n3622), .SI(n9544), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[1][114] ), .QN(n9543));
   SDFFARX1 \key_mem_reg[2][114]  (.D(n3623), .SI(n9416), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[2][114] ), .QN(n9415));
   SDFFARX1 \key_mem_reg[3][114]  (.D(n3624), .SI(n9288), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[3][114] ), .QN(n9287));
   SDFFARX1 \key_mem_reg[4][114]  (.D(n3625), .SI(n9161), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[4][114] ), .QN(n9160));
   SDFFARX1 \key_mem_reg[5][114]  (.D(n3626), .SI(n9033), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[5][114] ), .QN(n9032));
   SDFFARX1 \key_mem_reg[6][114]  (.D(n3627), .SI(n8905), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[6][114] ), .QN(n8904));
   SDFFARX1 \key_mem_reg[7][114]  (.D(n3628), .SI(n8777), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[7][114] ), .QN(n8776));
   SDFFARX1 \key_mem_reg[8][114]  (.D(n3629), .SI(n8649), .SE(test_se), .CLK(clk), .RSTB(
          n7475), .Q(\key_mem[8][114] ), .QN(n8648));
   SDFFARX1 \key_mem_reg[9][114]  (.D(n3630), .SI(n8521), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[9][114] ), .QN(n8520));
   SDFFARX1 \key_mem_reg[10][114]  (.D(n3631), .SI(n8393), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[10][114] ), .QN(n8392));
   SDFFARX1 \key_mem_reg[11][114]  (.D(n3632), .SI(n8265), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[11][114] ), .QN(n8264));
   SDFFARX1 \key_mem_reg[12][114]  (.D(n3633), .SI(n8138), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[12][114] ), .QN(n8137));
   SDFFARX1 \key_mem_reg[13][114]  (.D(n3634), .SI(n8010), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[13][114] ), .QN(n8009));
   SDFFARX1 \key_mem_reg[14][114]  (.D(n3635), .SI(n7882), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[14][114] ), .QN(n7881));
   SDFFARX1 \prev_key1_reg_reg[113]  (.D(n5360), .SI(n7648), .SE(test_se), .CLK(clk), .
          RSTB(n7474), .Q(prev_key1_reg[113]), .QN(n7647));
   SDFFARX1 \prev_key0_reg_reg[113]  (.D(n5487), .SI(prev_key0_reg[112]), .SE(test_se), .
          CLK(clk), .RSTB(n7474), .Q(prev_key0_reg[113]), .QN(n2229));
   SDFFARX1 \key_mem_reg[0][113]  (.D(n3636), .SI(n9673), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[0][113] ), .QN(n9672));
   SDFFARX1 \key_mem_reg[1][113]  (.D(n3637), .SI(n9545), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[1][113] ), .QN(n9544));
   SDFFARX1 \key_mem_reg[2][113]  (.D(n3638), .SI(n9417), .SE(test_se), .CLK(clk), .RSTB(
          n7474), .Q(\key_mem[2][113] ), .QN(n9416));
   SDFFARX1 \key_mem_reg[3][113]  (.D(n3639), .SI(n9289), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7474), .Q(\key_mem[3][113] ), .QN(n9288));
   SDFFARX1 \key_mem_reg[4][113]  (.D(n3640), .SI(n9162), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[4][113] ), .QN(n9161));
   SDFFARX1 \key_mem_reg[5][113]  (.D(n3641), .SI(n9034), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[5][113] ), .QN(n9033));
   SDFFARX1 \key_mem_reg[6][113]  (.D(n3642), .SI(n8906), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[6][113] ), .QN(n8905));
   SDFFARX1 \key_mem_reg[7][113]  (.D(n3643), .SI(n8778), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[7][113] ), .QN(n8777));
   SDFFARX1 \key_mem_reg[8][113]  (.D(n3644), .SI(n8650), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[8][113] ), .QN(n8649));
   SDFFARX1 \key_mem_reg[9][113]  (.D(n3645), .SI(n8522), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[9][113] ), .QN(n8521));
   SDFFARX1 \key_mem_reg[10][113]  (.D(n3646), .SI(n8394), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[10][113] ), .QN(n8393));
   SDFFARX1 \key_mem_reg[11][113]  (.D(n3647), .SI(n8266), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[11][113] ), .QN(n8265));
   SDFFARX1 \key_mem_reg[12][113]  (.D(n3648), .SI(n8139), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[12][113] ), .QN(n8138));
   SDFFARX1 \key_mem_reg[13][113]  (.D(n3649), .SI(n8011), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[13][113] ), .QN(n8010));
   SDFFARX1 \key_mem_reg[14][113]  (.D(n3650), .SI(n7883), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(\key_mem[14][113] ), .QN(n7882));
   SDFFARX1 \prev_key1_reg_reg[112]  (.D(n5361), .SI(n2200), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7473), .Q(prev_key1_reg[112]), .QN(n7648));
   SDFFARX1 \prev_key0_reg_reg[112]  (.D(n5488), .SI(n7756), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(prev_key0_reg[112]), .QN(n2230));
   SDFFARX1 \key_mem_reg[0][112]  (.D(n3651), .SI(n9674), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[0][112] ), .QN(n9673));
   SDFFARX1 \key_mem_reg[1][112]  (.D(n3652), .SI(n9546), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[1][112] ), .QN(n9545));
   SDFFARX1 \key_mem_reg[2][112]  (.D(n3653), .SI(n9418), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[2][112] ), .QN(n9417));
   SDFFARX1 \key_mem_reg[3][112]  (.D(n3654), .SI(n9290), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[3][112] ), .QN(n9289));
   SDFFARX1 \key_mem_reg[4][112]  (.D(n3655), .SI(n9163), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[4][112] ), .QN(n9162));
   SDFFARX1 \key_mem_reg[5][112]  (.D(n3656), .SI(n9035), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[5][112] ), .QN(n9034));
   SDFFARX1 \key_mem_reg[6][112]  (.D(n3657), .SI(n8907), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[6][112] ), .QN(n8906));
   SDFFARX1 \key_mem_reg[7][112]  (.D(n3658), .SI(n8779), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[7][112] ), .QN(n8778));
   SDFFARX1 \key_mem_reg[8][112]  (.D(n3659), .SI(n8651), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[8][112] ), .QN(n8650));
   SDFFARX1 \key_mem_reg[9][112]  (.D(n3660), .SI(n8523), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[9][112] ), .QN(n8522));
   SDFFARX1 \key_mem_reg[10][112]  (.D(n3661), .SI(n8395), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7472), .Q(\key_mem[10][112] ), .QN(n8394));
   SDFFARX1 \key_mem_reg[11][112]  (.D(n3662), .SI(n8267), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[11][112] ), .QN(n8266));
   SDFFARX1 \key_mem_reg[12][112]  (.D(n3663), .SI(n8140), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[12][112] ), .QN(n8139));
   SDFFARX1 \key_mem_reg[13][112]  (.D(n3664), .SI(n8012), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[13][112] ), .QN(n8011));
   SDFFARX1 \key_mem_reg[14][112]  (.D(n3665), .SI(n7884), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[14][112] ), .QN(n7883));
   SDFFARX1 \prev_key1_reg_reg[111]  (.D(n5362), .SI(n7649), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(prev_key1_reg[111]), .QN(n2200));
   SDFFARX1 \prev_key0_reg_reg[111]  (.D(n5489), .SI(n7757), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(prev_key0_reg[111]), .QN(n7756));
   SDFFARX1 \key_mem_reg[0][111]  (.D(n3666), .SI(n9675), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[0][111] ), .QN(n9674));
   SDFFARX1 \key_mem_reg[1][111]  (.D(n3667), .SI(n9547), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[1][111] ), .QN(n9546));
   SDFFARX1 \key_mem_reg[2][111]  (.D(n3668), .SI(n9419), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[2][111] ), .QN(n9418));
   SDFFARX1 \key_mem_reg[3][111]  (.D(n3669), .SI(n9291), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[3][111] ), .QN(n9290));
   SDFFARX1 \key_mem_reg[4][111]  (.D(n3670), .SI(n9164), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[4][111] ), .QN(n9163));
   SDFFARX1 \key_mem_reg[5][111]  (.D(n3671), .SI(n9036), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7471), .Q(\key_mem[5][111] ), .QN(n9035));
   SDFFARX1 \key_mem_reg[6][111]  (.D(n3672), .SI(n8908), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[6][111] ), .QN(n8907));
   SDFFARX1 \key_mem_reg[7][111]  (.D(n3673), .SI(n8780), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[7][111] ), .QN(n8779));
   SDFFARX1 \key_mem_reg[8][111]  (.D(n3674), .SI(n8652), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[8][111] ), .QN(n8651));
   SDFFARX1 \key_mem_reg[9][111]  (.D(n3675), .SI(n8524), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[9][111] ), .QN(n8523));
   SDFFARX1 \key_mem_reg[10][111]  (.D(n3676), .SI(n8396), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[10][111] ), .QN(n8395));
   SDFFARX1 \key_mem_reg[11][111]  (.D(n3677), .SI(n8268), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[11][111] ), .QN(n8267));
   SDFFARX1 \key_mem_reg[12][111]  (.D(n3678), .SI(n8141), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[12][111] ), .QN(n8140));
   SDFFARX1 \key_mem_reg[13][111]  (.D(n3679), .SI(n8013), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[13][111] ), .QN(n8012));
   SDFFARX1 \key_mem_reg[14][111]  (.D(n3680), .SI(n7885), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[14][111] ), .QN(n7884));
   SDFFARX1 \prev_key1_reg_reg[110]  (.D(n5363), .SI(n2198), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(prev_key1_reg[110]), .QN(n7649));
   SDFFARX1 \prev_key0_reg_reg[110]  (.D(n5490), .SI(n7758), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(prev_key0_reg[110]), .QN(n7757));
   SDFFARX1 \key_mem_reg[0][110]  (.D(n3681), .SI(n9676), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7470), .Q(\key_mem[0][110] ), .QN(n9675));
   SDFFARX1 \key_mem_reg[2][110]  (.D(n3683), .SI(n9420), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[2][110] ), .QN(n9419));
   SDFFARX1 \key_mem_reg[3][110]  (.D(n3684), .SI(n9292), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[3][110] ), .QN(n9291));
   SDFFARX1 \key_mem_reg[4][110]  (.D(n3685), .SI(n9165), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[4][110] ), .QN(n9164));
   SDFFARX1 \key_mem_reg[5][110]  (.D(n3686), .SI(n9037), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[5][110] ), .QN(n9036));
   SDFFARX1 \key_mem_reg[6][110]  (.D(n3687), .SI(n8909), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[6][110] ), .QN(n8908));
   SDFFARX1 \key_mem_reg[7][110]  (.D(n3688), .SI(n8781), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[7][110] ), .QN(n8780));
   SDFFARX1 \key_mem_reg[8][110]  (.D(n3689), .SI(n8653), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[8][110] ), .QN(n8652));
   SDFFARX1 \key_mem_reg[9][110]  (.D(n3690), .SI(n8525), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[9][110] ), .QN(n8524));
   SDFFARX1 \key_mem_reg[10][110]  (.D(n3691), .SI(n8397), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[10][110] ), .QN(n8396));
   SDFFARX1 \key_mem_reg[11][110]  (.D(n3692), .SI(n8269), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[11][110] ), .QN(n8268));
   SDFFARX1 \key_mem_reg[12][110]  (.D(n3693), .SI(n8142), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7469), .Q(\key_mem[12][110] ), .QN(n8141));
   SDFFARX1 \key_mem_reg[13][110]  (.D(n3694), .SI(n8014), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[13][110] ), .QN(n8013));
   SDFFARX1 \key_mem_reg[14][110]  (.D(n3695), .SI(n7886), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[14][110] ), .QN(n7885));
   SDFFARX1 \prev_key1_reg_reg[109]  (.D(n5364), .SI(n7650), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(prev_key1_reg[109]), .QN(n2198));
   SDFFARX1 \prev_key0_reg_reg[109]  (.D(n5491), .SI(n7759), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(prev_key0_reg[109]), .QN(n7758));
   SDFFARX1 \key_mem_reg[0][109]  (.D(n3696), .SI(n9677), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[0][109] ), .QN(n9676));
   SDFFARX1 \key_mem_reg[1][109]  (.D(n3697), .SI(n9549), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[1][109] ), .QN(n9548));
   SDFFARX1 \key_mem_reg[2][109]  (.D(n3698), .SI(n9421), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[2][109] ), .QN(n9420));
   SDFFARX1 \key_mem_reg[3][109]  (.D(n3699), .SI(n9293), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[3][109] ), .QN(n9292));
   SDFFARX1 \key_mem_reg[4][109]  (.D(n3700), .SI(n9166), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[4][109] ), .QN(n9165));
   SDFFARX1 \key_mem_reg[5][109]  (.D(n3701), .SI(n9038), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[5][109] ), .QN(n9037));
   SDFFARX1 \key_mem_reg[6][109]  (.D(n3702), .SI(n8910), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[6][109] ), .QN(n8909));
   SDFFARX1 \key_mem_reg[7][109]  (.D(n3703), .SI(n8782), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7468), .Q(\key_mem[7][109] ), .QN(n8781));
   SDFFARX1 \key_mem_reg[8][109]  (.D(n3704), .SI(n8654), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[8][109] ), .QN(n8653));
   SDFFARX1 \key_mem_reg[9][109]  (.D(n3705), .SI(n8526), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[9][109] ), .QN(n8525));
   SDFFARX1 \key_mem_reg[10][109]  (.D(n3706), .SI(n8398), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[10][109] ), .QN(n8397));
   SDFFARX1 \key_mem_reg[11][109]  (.D(n3707), .SI(n8270), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[11][109] ), .QN(n8269));
   SDFFARX1 \key_mem_reg[12][109]  (.D(n3708), .SI(n8143), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[12][109] ), .QN(n8142));
   SDFFARX1 \key_mem_reg[13][109]  (.D(n3709), .SI(n8015), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[13][109] ), .QN(n8014));
   SDFFARX1 \key_mem_reg[14][109]  (.D(n3710), .SI(n7887), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[14][109] ), .QN(n7886));
   SDFFARX1 \prev_key1_reg_reg[108]  (.D(n5365), .SI(n7651), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(prev_key1_reg[108]), .QN(n7650));
   SDFFARX1 \prev_key0_reg_reg[108]  (.D(n5492), .SI(n7760), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(prev_key0_reg[108]), .QN(n7759));
   SDFFARX1 \key_mem_reg[0][108]  (.D(n3711), .SI(n9678), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[0][108] ), .QN(n9677));
   SDFFARX1 \key_mem_reg[1][108]  (.D(n3712), .SI(n9550), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[1][108] ), .QN(n9549));
   SDFFARX1 \key_mem_reg[2][108]  (.D(n3713), .SI(n9422), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7467), .Q(\key_mem[2][108] ), .QN(n9421));
   SDFFARX1 \key_mem_reg[3][108]  (.D(n3714), .SI(n9294), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[3][108] ), .QN(n9293));
   SDFFARX1 \key_mem_reg[4][108]  (.D(n3715), .SI(n9167), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[4][108] ), .QN(n9166));
   SDFFARX1 \key_mem_reg[5][108]  (.D(n3716), .SI(n9039), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[5][108] ), .QN(n9038));
   SDFFARX1 \key_mem_reg[6][108]  (.D(n3717), .SI(n8911), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[6][108] ), .QN(n8910));
   SDFFARX1 \key_mem_reg[7][108]  (.D(n3718), .SI(n8783), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[7][108] ), .QN(n8782));
   SDFFARX1 \key_mem_reg[8][108]  (.D(n3719), .SI(n8655), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[8][108] ), .QN(n8654));
   SDFFARX1 \key_mem_reg[9][108]  (.D(n3720), .SI(n8527), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[9][108] ), .QN(n8526));
   SDFFARX1 \key_mem_reg[10][108]  (.D(n3721), .SI(n8399), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[10][108] ), .QN(n8398));
   SDFFARX1 \key_mem_reg[11][108]  (.D(n3722), .SI(n8271), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[11][108] ), .QN(n8270));
   SDFFARX1 \key_mem_reg[12][108]  (.D(n3723), .SI(n8144), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[12][108] ), .QN(n8143));
   SDFFARX1 \key_mem_reg[13][108]  (.D(n3724), .SI(n8016), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[13][108] ), .QN(n8015));
   SDFFARX1 \key_mem_reg[14][108]  (.D(n3725), .SI(n7888), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7466), .Q(\key_mem[14][108] ), .QN(n7887));
   SDFFARX1 \prev_key1_reg_reg[107]  (.D(n5366), .SI(n2202), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(prev_key1_reg[107]), .QN(n7651));
   SDFFARX1 \prev_key0_reg_reg[107]  (.D(n5493), .SI(n7761), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(prev_key0_reg[107]), .QN(n7760));
   SDFFARX1 \key_mem_reg[0][107]  (.D(n3726), .SI(n9679), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[0][107] ), .QN(n9678));
   SDFFARX1 \key_mem_reg[1][107]  (.D(n3727), .SI(n9551), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[1][107] ), .QN(n9550));
   SDFFARX1 \key_mem_reg[2][107]  (.D(n3728), .SI(n9423), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[2][107] ), .QN(n9422));
   SDFFARX1 \key_mem_reg[3][107]  (.D(n3729), .SI(n9295), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[3][107] ), .QN(n9294));
   SDFFARX1 \key_mem_reg[4][107]  (.D(n3730), .SI(n9168), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[4][107] ), .QN(n9167));
   SDFFARX1 \key_mem_reg[5][107]  (.D(n3731), .SI(n9040), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[5][107] ), .QN(n9039));
   SDFFARX1 \key_mem_reg[6][107]  (.D(n3732), .SI(n8912), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[6][107] ), .QN(n8911));
   SDFFARX1 \key_mem_reg[7][107]  (.D(n3733), .SI(n8784), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[7][107] ), .QN(n8783));
   SDFFARX1 \key_mem_reg[8][107]  (.D(n3734), .SI(n8656), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[8][107] ), .QN(n8655));
   SDFFARX1 \key_mem_reg[9][107]  (.D(n3735), .SI(n8528), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7465), .Q(\key_mem[9][107] ), .QN(n8527));
   SDFFARX1 \key_mem_reg[10][107]  (.D(n3736), .SI(n8400), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[10][107] ), .QN(n8399));
   SDFFARX1 \key_mem_reg[11][107]  (.D(n3737), .SI(n8272), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[11][107] ), .QN(n8271));
   SDFFARX1 \key_mem_reg[12][107]  (.D(n3738), .SI(n8145), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[12][107] ), .QN(n8144));
   SDFFARX1 \key_mem_reg[13][107]  (.D(n3739), .SI(n8017), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[13][107] ), .QN(n8016));
   SDFFARX1 \key_mem_reg[14][107]  (.D(n3740), .SI(n7889), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[14][107] ), .QN(n7888));
   SDFFARX1 \prev_key1_reg_reg[106]  (.D(n5367), .SI(n7652), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(prev_key1_reg[106]), .QN(n2202));
   SDFFARX1 \prev_key0_reg_reg[106]  (.D(n5494), .SI(n7762), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(prev_key0_reg[106]), .QN(n7761));
   SDFFARX1 \key_mem_reg[0][106]  (.D(n3741), .SI(n9680), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[0][106] ), .QN(n9679));
   SDFFARX1 \key_mem_reg[1][106]  (.D(n3742), .SI(n9552), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[1][106] ), .QN(n9551));
   SDFFARX1 \key_mem_reg[2][106]  (.D(n3743), .SI(n9424), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[2][106] ), .QN(n9423));
   SDFFARX1 \key_mem_reg[3][106]  (.D(n3744), .SI(n9296), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[3][106] ), .QN(n9295));
   SDFFARX1 \key_mem_reg[4][106]  (.D(n3745), .SI(n9169), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7464), .Q(\key_mem[4][106] ), .QN(n9168));
   SDFFARX1 \key_mem_reg[5][106]  (.D(n3746), .SI(n9041), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[5][106] ), .QN(n9040));
   SDFFARX1 \key_mem_reg[6][106]  (.D(n3747), .SI(n8913), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[6][106] ), .QN(n8912));
   SDFFARX1 \key_mem_reg[7][106]  (.D(n3748), .SI(n8785), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[7][106] ), .QN(n8784));
   SDFFARX1 \key_mem_reg[8][106]  (.D(n3749), .SI(n8657), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[8][106] ), .QN(n8656));
   SDFFARX1 \key_mem_reg[9][106]  (.D(n3750), .SI(n8529), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[9][106] ), .QN(n8528));
   SDFFARX1 \key_mem_reg[10][106]  (.D(n3751), .SI(n8401), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[10][106] ), .QN(n8400));
   SDFFARX1 \key_mem_reg[11][106]  (.D(n3752), .SI(n8273), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[11][106] ), .QN(n8272));
   SDFFARX1 \key_mem_reg[12][106]  (.D(n3753), .SI(n8146), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[12][106] ), .QN(n8145));
   SDFFARX1 \key_mem_reg[13][106]  (.D(n3754), .SI(n8018), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[13][106] ), .QN(n8017));
   SDFFARX1 \key_mem_reg[14][106]  (.D(n3755), .SI(n7890), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(\key_mem[14][106] ), .QN(n7889));
   SDFFARX1 \prev_key1_reg_reg[105]  (.D(n5368), .SI(n7653), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(prev_key1_reg[105]), .QN(n7652));
   SDFFARX1 \prev_key0_reg_reg[105]  (.D(n5495), .SI(n7763), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7463), .Q(prev_key0_reg[105]), .QN(n7762));
   SDFFARX1 \key_mem_reg[0][105]  (.D(n3756), .SI(n9681), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[0][105] ), .QN(n9680));
   SDFFARX1 \key_mem_reg[1][105]  (.D(n3757), .SI(n9553), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[1][105] ), .QN(n9552));
   SDFFARX1 \key_mem_reg[2][105]  (.D(n3758), .SI(n9425), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[2][105] ), .QN(n9424));
   SDFFARX1 \key_mem_reg[3][105]  (.D(n3759), .SI(n9297), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[3][105] ), .QN(n9296));
   SDFFARX1 \key_mem_reg[4][105]  (.D(n3760), .SI(n9170), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[4][105] ), .QN(n9169));
   SDFFARX1 \key_mem_reg[5][105]  (.D(n3761), .SI(n9042), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[5][105] ), .QN(n9041));
   SDFFARX1 \key_mem_reg[6][105]  (.D(n3762), .SI(n8914), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[6][105] ), .QN(n8913));
   SDFFARX1 \key_mem_reg[7][105]  (.D(n3763), .SI(n8786), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[7][105] ), .QN(n8785));
   SDFFARX1 \key_mem_reg[8][105]  (.D(n3764), .SI(n8658), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[8][105] ), .QN(n8657));
   SDFFARX1 \key_mem_reg[9][105]  (.D(n3765), .SI(n8530), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[9][105] ), .QN(n8529));
   SDFFARX1 \key_mem_reg[10][105]  (.D(n3766), .SI(n8402), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[10][105] ), .QN(n8401));
   SDFFARX1 \key_mem_reg[11][105]  (.D(n3767), .SI(n8274), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7462), .Q(\key_mem[11][105] ), .QN(n8273));
   SDFFARX1 \key_mem_reg[12][105]  (.D(n3768), .SI(n8147), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[12][105] ), .QN(n8146));
   SDFFARX1 \key_mem_reg[13][105]  (.D(n3769), .SI(n8019), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[13][105] ), .QN(n8018));
   SDFFARX1 \key_mem_reg[14][105]  (.D(n3770), .SI(n7891), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[14][105] ), .QN(n7890));
   SDFFARX1 \prev_key1_reg_reg[104]  (.D(n5369), .SI(n7654), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(prev_key1_reg[104]), .QN(n7653));
   SDFFARX1 \prev_key0_reg_reg[104]  (.D(n5496), .SI(n7764), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(prev_key0_reg[104]), .QN(n7763));
   SDFFARX1 \key_mem_reg[0][104]  (.D(n3771), .SI(n9682), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[0][104] ), .QN(n9681));
   SDFFARX1 \key_mem_reg[1][104]  (.D(n3772), .SI(n9554), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[1][104] ), .QN(n9553));
   SDFFARX1 \key_mem_reg[2][104]  (.D(n3773), .SI(n9426), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[2][104] ), .QN(n9425));
   SDFFARX1 \key_mem_reg[3][104]  (.D(n3774), .SI(n9298), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[3][104] ), .QN(n9297));
   SDFFARX1 \key_mem_reg[4][104]  (.D(n3775), .SI(n9171), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[4][104] ), .QN(n9170));
   SDFFARX1 \key_mem_reg[5][104]  (.D(n3776), .SI(n9043), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[5][104] ), .QN(n9042));
   SDFFARX1 \key_mem_reg[6][104]  (.D(n3777), .SI(n8915), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7461), .Q(\key_mem[6][104] ), .QN(n8914));
   SDFFARX1 \key_mem_reg[7][104]  (.D(n3778), .SI(n8787), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[7][104] ), .QN(n8786));
   SDFFARX1 \key_mem_reg[8][104]  (.D(n3779), .SI(n8659), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[8][104] ), .QN(n8658));
   SDFFARX1 \key_mem_reg[9][104]  (.D(n3780), .SI(n8531), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[9][104] ), .QN(n8530));
   SDFFARX1 \key_mem_reg[10][104]  (.D(n3781), .SI(n8403), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[10][104] ), .QN(n8402));
   SDFFARX1 \key_mem_reg[11][104]  (.D(n3782), .SI(n8275), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[11][104] ), .QN(n8274));
   SDFFARX1 \key_mem_reg[12][104]  (.D(n3783), .SI(n8148), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[12][104] ), .QN(n8147));
   SDFFARX1 \key_mem_reg[13][104]  (.D(n3784), .SI(n8020), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[13][104] ), .QN(n8019));
   SDFFARX1 \key_mem_reg[14][104]  (.D(n3785), .SI(n7892), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[14][104] ), .QN(n7891));
   SDFFARX1 \prev_key1_reg_reg[103]  (.D(n5370), .SI(n7655), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(prev_key1_reg[103]), .QN(n7654));
   SDFFARX1 \prev_key0_reg_reg[103]  (.D(n5497), .SI(n7765), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(prev_key0_reg[103]), .QN(n7764));
   SDFFARX1 \key_mem_reg[0][103]  (.D(n3786), .SI(n9683), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[0][103] ), .QN(n9682));
   SDFFARX1 \key_mem_reg[1][103]  (.D(n3787), .SI(n9555), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7460), .Q(\key_mem[1][103] ), .QN(n9554));
   SDFFARX1 \key_mem_reg[2][103]  (.D(n3788), .SI(n9427), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[2][103] ), .QN(n9426));
   SDFFARX1 \key_mem_reg[3][103]  (.D(n3789), .SI(n9299), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[3][103] ), .QN(n9298));
   SDFFARX1 \key_mem_reg[4][103]  (.D(n3790), .SI(n9172), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[4][103] ), .QN(n9171));
   SDFFARX1 \key_mem_reg[5][103]  (.D(n3791), .SI(n9044), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[5][103] ), .QN(n9043));
   SDFFARX1 \key_mem_reg[6][103]  (.D(n3792), .SI(n8916), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[6][103] ), .QN(n8915));
   SDFFARX1 \key_mem_reg[7][103]  (.D(n3793), .SI(n8788), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[7][103] ), .QN(n8787));
   SDFFARX1 \key_mem_reg[8][103]  (.D(n3794), .SI(n8660), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[8][103] ), .QN(n8659));
   SDFFARX1 \key_mem_reg[9][103]  (.D(n3795), .SI(n8532), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[9][103] ), .QN(n8531));
   SDFFARX1 \key_mem_reg[10][103]  (.D(n3796), .SI(n8404), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[10][103] ), .QN(n8403));
   SDFFARX1 \key_mem_reg[11][103]  (.D(n3797), .SI(n8276), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[11][103] ), .QN(n8275));
   SDFFARX1 \key_mem_reg[12][103]  (.D(n3798), .SI(n8149), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[12][103] ), .QN(n8148));
   SDFFARX1 \key_mem_reg[13][103]  (.D(n3799), .SI(n8021), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7459), .Q(\key_mem[13][103] ), .QN(n8020));
   SDFFARX1 \key_mem_reg[14][103]  (.D(n3800), .SI(n7893), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[14][103] ), .QN(n7892));
   SDFFARX1 \prev_key1_reg_reg[102]  (.D(n5371), .SI(n7656), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(prev_key1_reg[102]), .QN(n7655));
   SDFFARX1 \prev_key0_reg_reg[102]  (.D(n5498), .SI(n7766), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(prev_key0_reg[102]), .QN(n7765));
   SDFFARX1 \key_mem_reg[0][102]  (.D(n3801), .SI(n9684), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[0][102] ), .QN(n9683));
   SDFFARX1 \key_mem_reg[1][102]  (.D(n3802), .SI(n9556), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[1][102] ), .QN(n9555));
   SDFFARX1 \key_mem_reg[2][102]  (.D(n3803), .SI(n9428), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[2][102] ), .QN(n9427));
   SDFFARX1 \key_mem_reg[3][102]  (.D(n3804), .SI(n9300), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[3][102] ), .QN(n9299));
   SDFFARX1 \key_mem_reg[4][102]  (.D(n3805), .SI(n9173), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[4][102] ), .QN(n9172));
   SDFFARX1 \key_mem_reg[5][102]  (.D(n3806), .SI(n9045), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[5][102] ), .QN(n9044));
   SDFFARX1 \key_mem_reg[6][102]  (.D(n3807), .SI(n8917), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[6][102] ), .QN(n8916));
   SDFFARX1 \key_mem_reg[7][102]  (.D(n3808), .SI(n8789), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[7][102] ), .QN(n8788));
   SDFFARX1 \key_mem_reg[8][102]  (.D(n3809), .SI(n8661), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7458), .Q(\key_mem[8][102] ), .QN(n8660));
   SDFFARX1 \key_mem_reg[9][102]  (.D(n3810), .SI(n8533), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[9][102] ), .QN(n8532));
   SDFFARX1 \key_mem_reg[10][102]  (.D(n3811), .SI(n8405), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[10][102] ), .QN(n8404));
   SDFFARX1 \key_mem_reg[11][102]  (.D(n3812), .SI(n8277), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[11][102] ), .QN(n8276));
   SDFFARX1 \key_mem_reg[12][102]  (.D(n3813), .SI(n8150), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[12][102] ), .QN(n8149));
   SDFFARX1 \key_mem_reg[13][102]  (.D(n3814), .SI(n8022), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[13][102] ), .QN(n8021));
   SDFFARX1 \key_mem_reg[14][102]  (.D(n3815), .SI(n7894), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[14][102] ), .QN(n7893));
   SDFFARX1 \prev_key1_reg_reg[101]  (.D(n5372), .SI(n7657), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(prev_key1_reg[101]), .QN(n7656));
   SDFFARX1 \prev_key0_reg_reg[101]  (.D(n5499), .SI(n7767), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(prev_key0_reg[101]), .QN(n7766));
   SDFFARX1 \key_mem_reg[0][101]  (.D(n3816), .SI(n9685), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[0][101] ), .QN(n9684));
   SDFFARX1 \key_mem_reg[1][101]  (.D(n3817), .SI(n9557), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[1][101] ), .QN(n9556));
   SDFFARX1 \key_mem_reg[2][101]  (.D(n3818), .SI(n9429), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[2][101] ), .QN(n9428));
   SDFFARX1 \key_mem_reg[3][101]  (.D(n3819), .SI(n9301), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7457), .Q(\key_mem[3][101] ), .QN(n9300));
   SDFFARX1 \key_mem_reg[4][101]  (.D(n3820), .SI(n9174), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[4][101] ), .QN(n9173));
   SDFFARX1 \key_mem_reg[5][101]  (.D(n3821), .SI(n9046), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[5][101] ), .QN(n9045));
   SDFFARX1 \key_mem_reg[6][101]  (.D(n3822), .SI(n8918), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[6][101] ), .QN(n8917));
   SDFFARX1 \key_mem_reg[7][101]  (.D(n3823), .SI(n8790), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[7][101] ), .QN(n8789));
   SDFFARX1 \key_mem_reg[8][101]  (.D(n3824), .SI(n8662), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[8][101] ), .QN(n8661));
   SDFFARX1 \key_mem_reg[9][101]  (.D(n3825), .SI(n8534), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[9][101] ), .QN(n8533));
   SDFFARX1 \key_mem_reg[10][101]  (.D(n3826), .SI(n8406), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[10][101] ), .QN(n8405));
   SDFFARX1 \key_mem_reg[11][101]  (.D(n3827), .SI(n8278), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[11][101] ), .QN(n8277));
   SDFFARX1 \key_mem_reg[12][101]  (.D(n3828), .SI(n8151), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[12][101] ), .QN(n8150));
   SDFFARX1 \key_mem_reg[13][101]  (.D(n3829), .SI(n8023), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[13][101] ), .QN(n8022));
   SDFFARX1 \key_mem_reg[14][101]  (.D(n3830), .SI(n7895), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(\key_mem[14][101] ), .QN(n7894));
   SDFFARX1 \prev_key1_reg_reg[100]  (.D(n5373), .SI(n7658), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7456), .Q(prev_key1_reg[100]), .QN(n7657));
   SDFFARX1 \prev_key0_reg_reg[100]  (.D(n5500), .SI(n7768), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(prev_key0_reg[100]), .QN(n7767));
   SDFFARX1 \key_mem_reg[0][100]  (.D(n3831), .SI(n9686), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[0][100] ), .QN(n9685));
   SDFFARX1 \key_mem_reg[1][100]  (.D(n3832), .SI(n9558), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[1][100] ), .QN(n9557));
   SDFFARX1 \key_mem_reg[2][100]  (.D(n3833), .SI(n9430), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[2][100] ), .QN(n9429));
   SDFFARX1 \key_mem_reg[3][100]  (.D(n3834), .SI(n9302), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[3][100] ), .QN(n9301));
   SDFFARX1 \key_mem_reg[4][100]  (.D(n3835), .SI(n9175), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[4][100] ), .QN(n9174));
   SDFFARX1 \key_mem_reg[5][100]  (.D(n3836), .SI(n9047), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[5][100] ), .QN(n9046));
   SDFFARX1 \key_mem_reg[6][100]  (.D(n3837), .SI(n8919), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[6][100] ), .QN(n8918));
   SDFFARX1 \key_mem_reg[7][100]  (.D(n3838), .SI(n8791), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[7][100] ), .QN(n8790));
   SDFFARX1 \key_mem_reg[8][100]  (.D(n3839), .SI(n8663), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[8][100] ), .QN(n8662));
   SDFFARX1 \key_mem_reg[9][100]  (.D(n3840), .SI(n8535), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[9][100] ), .QN(n8534));
   SDFFARX1 \key_mem_reg[10][100]  (.D(n3841), .SI(n8407), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7455), .Q(\key_mem[10][100] ), .QN(n8406));
   SDFFARX1 \key_mem_reg[11][100]  (.D(n3842), .SI(n8279), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[11][100] ), .QN(n8278));
   SDFFARX1 \key_mem_reg[12][100]  (.D(n3843), .SI(n8152), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[12][100] ), .QN(n8151));
   SDFFARX1 \key_mem_reg[13][100]  (.D(n3844), .SI(n8024), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[13][100] ), .QN(n8023));
   SDFFARX1 \key_mem_reg[14][100]  (.D(n3845), .SI(n7896), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[14][100] ), .QN(n7895));
   SDFFARX1 \prev_key1_reg_reg[99]  (.D(n5374), .SI(n7659), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(prev_key1_reg[99]), .QN(n7658));
   SDFFARX1 \prev_key0_reg_reg[99]  (.D(n5501), .SI(n7769), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(prev_key0_reg[99]), .QN(n7768));
   SDFFARX1 \key_mem_reg[0][99]  (.D(n3846), .SI(n9687), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[0][99] ), .QN(n9686));
   SDFFARX1 \key_mem_reg[1][99]  (.D(n3847), .SI(n9559), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[1][99] ), .QN(n9558));
   SDFFARX1 \key_mem_reg[2][99]  (.D(n3848), .SI(n9431), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[2][99] ), .QN(n9430));
   SDFFARX1 \key_mem_reg[3][99]  (.D(n3849), .SI(n9303), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[3][99] ), .QN(n9302));
   SDFFARX1 \key_mem_reg[4][99]  (.D(n3850), .SI(n9176), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[4][99] ), .QN(n9175));
   SDFFARX1 \key_mem_reg[5][99]  (.D(n3851), .SI(n9048), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7454), .Q(\key_mem[5][99] ), .QN(n9047));
   SDFFARX1 \key_mem_reg[6][99]  (.D(n3852), .SI(n8920), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[6][99] ), .QN(n8919));
   SDFFARX1 \key_mem_reg[7][99]  (.D(n3853), .SI(n8792), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[7][99] ), .QN(n8791));
   SDFFARX1 \key_mem_reg[8][99]  (.D(n3854), .SI(n8664), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[8][99] ), .QN(n8663));
   SDFFARX1 \key_mem_reg[9][99]  (.D(n3855), .SI(n8536), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[9][99] ), .QN(n8535));
   SDFFARX1 \key_mem_reg[10][99]  (.D(n3856), .SI(n8408), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[10][99] ), .QN(n8407));
   SDFFARX1 \key_mem_reg[11][99]  (.D(n3857), .SI(n8280), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[11][99] ), .QN(n8279));
   SDFFARX1 \key_mem_reg[12][99]  (.D(n3858), .SI(n8153), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[12][99] ), .QN(n8152));
   SDFFARX1 \key_mem_reg[13][99]  (.D(n3859), .SI(n8025), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[13][99] ), .QN(n8024));
   SDFFARX1 \key_mem_reg[14][99]  (.D(n3860), .SI(n7897), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[14][99] ), .QN(n7896));
   SDFFARX1 \prev_key1_reg_reg[98]  (.D(n5375), .SI(n7660), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(prev_key1_reg[98]), .QN(n7659));
   SDFFARX1 \prev_key0_reg_reg[98]  (.D(n5502), .SI(n7770), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(prev_key0_reg[98]), .QN(n7769));
   SDFFARX1 \key_mem_reg[0][98]  (.D(n3861), .SI(n9688), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7453), .Q(\key_mem[0][98] ), .QN(n9687));
   SDFFARX1 \key_mem_reg[1][98]  (.D(n3862), .SI(n9560), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7452), .Q(\key_mem[1][98] ), .QN(n9559));
   SDFFARX1 \key_mem_reg[2][98]  (.D(n3863), .SI(n9432), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7452), .Q(\key_mem[2][98] ), .QN(n9431));
   SDFFARX1 \key_mem_reg[3][98]  (.D(n3864), .SI(n9304), .SE(test_se_buf_net0), .CLK(
          clk_buf_net0), .RSTB(n7452), .Q(\key_mem[3][98] ), .QN(n9303));
   SDFFARX1 \key_mem_reg[4][98]  (.D(n3865), .SI(n9177), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[4][98] ), .QN(n9176));
   SDFFARX1 \key_mem_reg[5][98]  (.D(n3866), .SI(n9049), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[5][98] ), .QN(n9048));
   SDFFARX1 \key_mem_reg[6][98]  (.D(n3867), .SI(n8921), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[6][98] ), .QN(n8920));
   SDFFARX1 \key_mem_reg[7][98]  (.D(n3868), .SI(n8793), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[7][98] ), .QN(n8792));
   SDFFARX1 \key_mem_reg[8][98]  (.D(n3869), .SI(n8665), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[8][98] ), .QN(n8664));
   SDFFARX1 \key_mem_reg[9][98]  (.D(n3870), .SI(n8537), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[9][98] ), .QN(n8536));
   SDFFARX1 \key_mem_reg[10][98]  (.D(n3871), .SI(n8409), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[10][98] ), .QN(n8408));
   SDFFARX1 \key_mem_reg[11][98]  (.D(n3872), .SI(n8281), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[11][98] ), .QN(n8280));
   SDFFARX1 \key_mem_reg[12][98]  (.D(n3873), .SI(n8154), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7452), .Q(\key_mem[12][98] ), .QN(n8153));
   SDFFARX1 \key_mem_reg[13][98]  (.D(n3874), .SI(n8026), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[13][98] ), .QN(n8025));
   SDFFARX1 \key_mem_reg[14][98]  (.D(n3875), .SI(n7898), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[14][98] ), .QN(n7897));
   SDFFARX1 \prev_key1_reg_reg[97]  (.D(n5376), .SI(n7661), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(prev_key1_reg[97]), .QN(n7660));
   SDFFARX1 \prev_key0_reg_reg[97]  (.D(n5503), .SI(n7771), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(prev_key0_reg[97]), .QN(n7770));
   SDFFARX1 \key_mem_reg[0][97]  (.D(n3876), .SI(n9689), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[0][97] ), .QN(n9688));
   SDFFARX1 \key_mem_reg[1][97]  (.D(n3877), .SI(n9561), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[1][97] ), .QN(n9560));
   SDFFARX1 \key_mem_reg[2][97]  (.D(n3878), .SI(n9433), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[2][97] ), .QN(n9432));
   SDFFARX1 \key_mem_reg[3][97]  (.D(n3879), .SI(n9305), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[3][97] ), .QN(n9304));
   SDFFARX1 \key_mem_reg[4][97]  (.D(n3880), .SI(n9178), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[4][97] ), .QN(n9177));
   SDFFARX1 \key_mem_reg[5][97]  (.D(n3881), .SI(n9050), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[5][97] ), .QN(n9049));
   SDFFARX1 \key_mem_reg[6][97]  (.D(n3882), .SI(n8922), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[6][97] ), .QN(n8921));
   SDFFARX1 \key_mem_reg[7][97]  (.D(n3883), .SI(n8794), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7451), .Q(\key_mem[7][97] ), .QN(n8793));
   SDFFARX1 \key_mem_reg[8][97]  (.D(n3884), .SI(n8666), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[8][97] ), .QN(n8665));
   SDFFARX1 \key_mem_reg[9][97]  (.D(n3885), .SI(n8538), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[9][97] ), .QN(n8537));
   SDFFARX1 \key_mem_reg[10][97]  (.D(n3886), .SI(n8410), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[10][97] ), .QN(n8409));
   SDFFARX1 \key_mem_reg[11][97]  (.D(n3887), .SI(n8282), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[11][97] ), .QN(n8281));
   SDFFARX1 \key_mem_reg[12][97]  (.D(n3888), .SI(n8155), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[12][97] ), .QN(n8154));
   SDFFARX1 \key_mem_reg[13][97]  (.D(n3889), .SI(n8027), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[13][97] ), .QN(n8026));
   SDFFARX1 \key_mem_reg[14][97]  (.D(n3890), .SI(n7899), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[14][97] ), .QN(n7898));
   SDFFARX1 \prev_key1_reg_reg[96]  (.D(n5377), .SI(n7662), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(prev_key1_reg[96]), .QN(n7661));
   SDFFARX1 \prev_key0_reg_reg[96]  (.D(n5504), .SI(n7772), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(prev_key0_reg[96]), .QN(n7771));
   SDFFARX1 \key_mem_reg[0][96]  (.D(n3891), .SI(n9690), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[0][96] ), .QN(n9689));
   SDFFARX1 \key_mem_reg[1][96]  (.D(n3892), .SI(n9562), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[1][96] ), .QN(n9561));
   SDFFARX1 \key_mem_reg[2][96]  (.D(n3893), .SI(n9434), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7450), .Q(\key_mem[2][96] ), .QN(n9433));
   SDFFARX1 \key_mem_reg[3][96]  (.D(n3894), .SI(n9306), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[3][96] ), .QN(n9305));
   SDFFARX1 \key_mem_reg[4][96]  (.D(n3895), .SI(n9179), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[4][96] ), .QN(n9178));
   SDFFARX1 \key_mem_reg[5][96]  (.D(n3896), .SI(n9051), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[5][96] ), .QN(n9050));
   SDFFARX1 \key_mem_reg[6][96]  (.D(n3897), .SI(n8923), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[6][96] ), .QN(n8922));
   SDFFARX1 \key_mem_reg[7][96]  (.D(n3898), .SI(n8795), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[7][96] ), .QN(n8794));
   SDFFARX1 \key_mem_reg[8][96]  (.D(n3899), .SI(n8667), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[8][96] ), .QN(n8666));
   SDFFARX1 \key_mem_reg[9][96]  (.D(n3900), .SI(n8539), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[9][96] ), .QN(n8538));
   SDFFARX1 \key_mem_reg[10][96]  (.D(n3901), .SI(n8411), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[10][96] ), .QN(n8410));
   SDFFARX1 \key_mem_reg[11][96]  (.D(n3902), .SI(n8283), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[11][96] ), .QN(n8282));
   SDFFARX1 \key_mem_reg[12][96]  (.D(n3903), .SI(n8156), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[12][96] ), .QN(n8155));
   SDFFARX1 \key_mem_reg[13][96]  (.D(n3904), .SI(n8028), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[13][96] ), .QN(n8027));
   SDFFARX1 \key_mem_reg[14][96]  (.D(n3905), .SI(n7900), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7449), .Q(\key_mem[14][96] ), .QN(n7899));
   SDFFARX1 \prev_key1_reg_reg[95]  (.D(n5378), .SI(n7663), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(prev_key1_reg[95]), .QN(n7662));
   SDFFARX1 \prev_key0_reg_reg[95]  (.D(n5505), .SI(n7773), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(prev_key0_reg[95]), .QN(n7772));
   SDFFARX1 \key_mem_reg[0][95]  (.D(n3906), .SI(n9691), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[0][95] ), .QN(n9690));
   SDFFARX1 \key_mem_reg[1][95]  (.D(n3907), .SI(n9563), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[1][95] ), .QN(n9562));
   SDFFARX1 \key_mem_reg[2][95]  (.D(n3908), .SI(n9435), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[2][95] ), .QN(n9434));
   SDFFARX1 \key_mem_reg[3][95]  (.D(n3909), .SI(n9307), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[3][95] ), .QN(n9306));
   SDFFARX1 \key_mem_reg[4][95]  (.D(n3910), .SI(n9180), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[4][95] ), .QN(n9179));
   SDFFARX1 \key_mem_reg[5][95]  (.D(n3911), .SI(n9052), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[5][95] ), .QN(n9051));
   SDFFARX1 \key_mem_reg[6][95]  (.D(n3912), .SI(n8924), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[6][95] ), .QN(n8923));
   SDFFARX1 \key_mem_reg[7][95]  (.D(n3913), .SI(n8796), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[7][95] ), .QN(n8795));
   SDFFARX1 \key_mem_reg[8][95]  (.D(n3914), .SI(n8668), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[8][95] ), .QN(n8667));
   SDFFARX1 \key_mem_reg[9][95]  (.D(n3915), .SI(n8540), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7448), .Q(\key_mem[9][95] ), .QN(n8539));
   SDFFARX1 \key_mem_reg[10][95]  (.D(n3916), .SI(n8412), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[10][95] ), .QN(n8411));
   SDFFARX1 \key_mem_reg[11][95]  (.D(n3917), .SI(n8284), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[11][95] ), .QN(n8283));
   SDFFARX1 \key_mem_reg[12][95]  (.D(n3918), .SI(n8157), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[12][95] ), .QN(n8156));
   SDFFARX1 \key_mem_reg[13][95]  (.D(n3919), .SI(n8029), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[13][95] ), .QN(n8028));
   SDFFARX1 \key_mem_reg[14][95]  (.D(n3920), .SI(n7901), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[14][95] ), .QN(n7900));
   SDFFARX1 \prev_key1_reg_reg[94]  (.D(n5379), .SI(n7664), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(prev_key1_reg[94]), .QN(n7663));
   SDFFARX1 \prev_key0_reg_reg[94]  (.D(n5506), .SI(n7774), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(prev_key0_reg[94]), .QN(n7773));
   SDFFARX1 \key_mem_reg[0][94]  (.D(n3921), .SI(n9692), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[0][94] ), .QN(n9691));
   SDFFARX1 \key_mem_reg[1][94]  (.D(n3922), .SI(n9564), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[1][94] ), .QN(n9563));
   SDFFARX1 \key_mem_reg[2][94]  (.D(n3923), .SI(n9436), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[2][94] ), .QN(n9435));
   SDFFARX1 \key_mem_reg[3][94]  (.D(n3924), .SI(n9308), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[3][94] ), .QN(n9307));
   SDFFARX1 \key_mem_reg[4][94]  (.D(n3925), .SI(n9181), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7447), .Q(\key_mem[4][94] ), .QN(n9180));
   SDFFARX1 \key_mem_reg[5][94]  (.D(n3926), .SI(n9053), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[5][94] ), .QN(n9052));
   SDFFARX1 \key_mem_reg[6][94]  (.D(n3927), .SI(n8925), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[6][94] ), .QN(n8924));
   SDFFARX1 \key_mem_reg[7][94]  (.D(n3928), .SI(n8797), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[7][94] ), .QN(n8796));
   SDFFARX1 \key_mem_reg[8][94]  (.D(n3929), .SI(n8669), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[8][94] ), .QN(n8668));
   SDFFARX1 \key_mem_reg[9][94]  (.D(n3930), .SI(n8541), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[9][94] ), .QN(n8540));
   SDFFARX1 \key_mem_reg[10][94]  (.D(n3931), .SI(n8413), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[10][94] ), .QN(n8412));
   SDFFARX1 \key_mem_reg[11][94]  (.D(n3932), .SI(n8285), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[11][94] ), .QN(n8284));
   SDFFARX1 \key_mem_reg[12][94]  (.D(n3933), .SI(n8158), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[12][94] ), .QN(n8157));
   SDFFARX1 \key_mem_reg[13][94]  (.D(n3934), .SI(n8030), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[13][94] ), .QN(n8029));
   SDFFARX1 \key_mem_reg[14][94]  (.D(n3935), .SI(n7902), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(\key_mem[14][94] ), .QN(n7901));
   SDFFARX1 \prev_key1_reg_reg[93]  (.D(n5380), .SI(n7665), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(prev_key1_reg[93]), .QN(n7664));
   SDFFARX1 \prev_key0_reg_reg[93]  (.D(n5507), .SI(n7775), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7446), .Q(prev_key0_reg[93]), .QN(n7774));
   SDFFARX1 \key_mem_reg[0][93]  (.D(n3936), .SI(n9693), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[0][93] ), .QN(n9692));
   SDFFARX1 \key_mem_reg[1][93]  (.D(n3937), .SI(n9565), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[1][93] ), .QN(n9564));
   SDFFARX1 \key_mem_reg[2][93]  (.D(n3938), .SI(n9437), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[2][93] ), .QN(n9436));
   SDFFARX1 \key_mem_reg[3][93]  (.D(n3939), .SI(n9309), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[3][93] ), .QN(n9308));
   SDFFARX1 \key_mem_reg[4][93]  (.D(n3940), .SI(n9182), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[4][93] ), .QN(n9181));
   SDFFARX1 \key_mem_reg[5][93]  (.D(n3941), .SI(n9054), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[5][93] ), .QN(n9053));
   SDFFARX1 \key_mem_reg[6][93]  (.D(n3942), .SI(n8926), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[6][93] ), .QN(n8925));
   SDFFARX1 \key_mem_reg[7][93]  (.D(n3943), .SI(n8798), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[7][93] ), .QN(n8797));
   SDFFARX1 \key_mem_reg[8][93]  (.D(n3944), .SI(n8670), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[8][93] ), .QN(n8669));
   SDFFARX1 \key_mem_reg[9][93]  (.D(n3945), .SI(n8542), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[9][93] ), .QN(n8541));
   SDFFARX1 \key_mem_reg[10][93]  (.D(n3946), .SI(n8414), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[10][93] ), .QN(n8413));
   SDFFARX1 \key_mem_reg[11][93]  (.D(n3947), .SI(n8286), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7445), .Q(\key_mem[11][93] ), .QN(n8285));
   SDFFARX1 \key_mem_reg[12][93]  (.D(n3948), .SI(n8159), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[12][93] ), .QN(n8158));
   SDFFARX1 \key_mem_reg[13][93]  (.D(n3949), .SI(n8031), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[13][93] ), .QN(n8030));
   SDFFARX1 \key_mem_reg[14][93]  (.D(n3950), .SI(n7903), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[14][93] ), .QN(n7902));
   SDFFARX1 \prev_key1_reg_reg[92]  (.D(n5381), .SI(n7666), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(prev_key1_reg[92]), .QN(n7665));
   SDFFARX1 \prev_key0_reg_reg[92]  (.D(n5508), .SI(n7776), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(prev_key0_reg[92]), .QN(n7775));
   SDFFARX1 \key_mem_reg[0][92]  (.D(n3951), .SI(n9694), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[0][92] ), .QN(n9693));
   SDFFARX1 \key_mem_reg[1][92]  (.D(n3952), .SI(n9566), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[1][92] ), .QN(n9565));
   SDFFARX1 \key_mem_reg[2][92]  (.D(n3953), .SI(n9438), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[2][92] ), .QN(n9437));
   SDFFARX1 \key_mem_reg[3][92]  (.D(n3954), .SI(n9310), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[3][92] ), .QN(n9309));
   SDFFARX1 \key_mem_reg[4][92]  (.D(n3955), .SI(n9183), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[4][92] ), .QN(n9182));
   SDFFARX1 \key_mem_reg[5][92]  (.D(n3956), .SI(n9055), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[5][92] ), .QN(n9054));
   SDFFARX1 \key_mem_reg[6][92]  (.D(n3957), .SI(n8927), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7444), .Q(\key_mem[6][92] ), .QN(n8926));
   SDFFARX1 \key_mem_reg[7][92]  (.D(n3958), .SI(n8799), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[7][92] ), .QN(n8798));
   SDFFARX1 \key_mem_reg[8][92]  (.D(n3959), .SI(n8671), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[8][92] ), .QN(n8670));
   SDFFARX1 \key_mem_reg[9][92]  (.D(n3960), .SI(n8543), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[9][92] ), .QN(n8542));
   SDFFARX1 \key_mem_reg[10][92]  (.D(n3961), .SI(n8415), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[10][92] ), .QN(n8414));
   SDFFARX1 \key_mem_reg[11][92]  (.D(n3962), .SI(n8287), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[11][92] ), .QN(n8286));
   SDFFARX1 \key_mem_reg[12][92]  (.D(n3963), .SI(n8160), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[12][92] ), .QN(n8159));
   SDFFARX1 \key_mem_reg[13][92]  (.D(n3964), .SI(n8032), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[13][92] ), .QN(n8031));
   SDFFARX1 \key_mem_reg[14][92]  (.D(n3965), .SI(n7904), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[14][92] ), .QN(n7903));
   SDFFARX1 \prev_key1_reg_reg[91]  (.D(n5382), .SI(n7667), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(prev_key1_reg[91]), .QN(n7666));
   SDFFARX1 \prev_key0_reg_reg[91]  (.D(n5509), .SI(n7777), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(prev_key0_reg[91]), .QN(n7776));
   SDFFARX1 \key_mem_reg[0][91]  (.D(n3966), .SI(n9695), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[0][91] ), .QN(n9694));
   SDFFARX1 \key_mem_reg[1][91]  (.D(n3967), .SI(n9567), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7443), .Q(\key_mem[1][91] ), .QN(n9566));
   SDFFARX1 \key_mem_reg[2][91]  (.D(n3968), .SI(n9439), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[2][91] ), .QN(n9438));
   SDFFARX1 \key_mem_reg[3][91]  (.D(n3969), .SI(n9311), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[3][91] ), .QN(n9310));
   SDFFARX1 \key_mem_reg[4][91]  (.D(n3970), .SI(n9184), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[4][91] ), .QN(n9183));
   SDFFARX1 \key_mem_reg[5][91]  (.D(n3971), .SI(n9056), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[5][91] ), .QN(n9055));
   SDFFARX1 \key_mem_reg[6][91]  (.D(n3972), .SI(n8928), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[6][91] ), .QN(n8927));
   SDFFARX1 \key_mem_reg[7][91]  (.D(n3973), .SI(n8800), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[7][91] ), .QN(n8799));
   SDFFARX1 \key_mem_reg[8][91]  (.D(n3974), .SI(n8672), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[8][91] ), .QN(n8671));
   SDFFARX1 \key_mem_reg[9][91]  (.D(n3975), .SI(n8544), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[9][91] ), .QN(n8543));
   SDFFARX1 \key_mem_reg[10][91]  (.D(n3976), .SI(n8416), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[10][91] ), .QN(n8415));
   SDFFARX1 \key_mem_reg[11][91]  (.D(n3977), .SI(n8288), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[11][91] ), .QN(n8287));
   SDFFARX1 \key_mem_reg[12][91]  (.D(n3978), .SI(n8161), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[12][91] ), .QN(n8160));
   SDFFARX1 \key_mem_reg[13][91]  (.D(n3979), .SI(n8033), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7442), .Q(\key_mem[13][91] ), .QN(n8032));
   SDFFARX1 \key_mem_reg[14][91]  (.D(n3980), .SI(n7905), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[14][91] ), .QN(n7904));
   SDFFARX1 \prev_key1_reg_reg[90]  (.D(n5383), .SI(n7668), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(prev_key1_reg[90]), .QN(n7667));
   SDFFARX1 \prev_key0_reg_reg[90]  (.D(n5510), .SI(n7778), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(prev_key0_reg[90]), .QN(n7777));
   SDFFARX1 \key_mem_reg[0][90]  (.D(n3981), .SI(n9696), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[0][90] ), .QN(n9695));
   SDFFARX1 \key_mem_reg[1][90]  (.D(n3982), .SI(n9568), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[1][90] ), .QN(n9567));
   SDFFARX1 \key_mem_reg[2][90]  (.D(n3983), .SI(n9440), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[2][90] ), .QN(n9439));
   SDFFARX1 \key_mem_reg[3][90]  (.D(n3984), .SI(n9312), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[3][90] ), .QN(n9311));
   SDFFARX1 \key_mem_reg[4][90]  (.D(n3985), .SI(n9185), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[4][90] ), .QN(n9184));
   SDFFARX1 \key_mem_reg[5][90]  (.D(n3986), .SI(n9057), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[5][90] ), .QN(n9056));
   SDFFARX1 \key_mem_reg[6][90]  (.D(n3987), .SI(n8929), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[6][90] ), .QN(n8928));
   SDFFARX1 \key_mem_reg[7][90]  (.D(n3988), .SI(n8801), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[7][90] ), .QN(n8800));
   SDFFARX1 \key_mem_reg[8][90]  (.D(n3989), .SI(n8673), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7441), .Q(\key_mem[8][90] ), .QN(n8672));
   SDFFARX1 \key_mem_reg[9][90]  (.D(n3990), .SI(n8545), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[9][90] ), .QN(n8544));
   SDFFARX1 \key_mem_reg[10][90]  (.D(n3991), .SI(n8417), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[10][90] ), .QN(n8416));
   SDFFARX1 \key_mem_reg[11][90]  (.D(n3992), .SI(n8289), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[11][90] ), .QN(n8288));
   SDFFARX1 \key_mem_reg[12][90]  (.D(n3993), .SI(n8162), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[12][90] ), .QN(n8161));
   SDFFARX1 \key_mem_reg[13][90]  (.D(n3994), .SI(n8034), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[13][90] ), .QN(n8033));
   SDFFARX1 \key_mem_reg[14][90]  (.D(n3995), .SI(n7906), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[14][90] ), .QN(n7905));
   SDFFARX1 \prev_key1_reg_reg[89]  (.D(n5384), .SI(n3), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(prev_key1_reg[89]), .QN(n7668));
   SDFFARX1 \prev_key0_reg_reg[89]  (.D(n5511), .SI(n7779), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(prev_key0_reg[89]), .QN(n7778));
   SDFFARX1 \key_mem_reg[0][89]  (.D(n3996), .SI(n9697), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[0][89] ), .QN(n9696));
   SDFFARX1 \key_mem_reg[1][89]  (.D(n3997), .SI(n9569), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[1][89] ), .QN(n9568));
   SDFFARX1 \key_mem_reg[2][89]  (.D(n3998), .SI(n9441), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[2][89] ), .QN(n9440));
   SDFFARX1 \key_mem_reg[3][89]  (.D(n3999), .SI(n9313), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7440), .Q(\key_mem[3][89] ), .QN(n9312));
   SDFFARX1 \key_mem_reg[4][89]  (.D(n4000), .SI(n9186), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[4][89] ), .QN(n9185));
   SDFFARX1 \key_mem_reg[5][89]  (.D(n4001), .SI(n9058), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[5][89] ), .QN(n9057));
   SDFFARX1 \key_mem_reg[6][89]  (.D(n4002), .SI(n8930), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[6][89] ), .QN(n8929));
   SDFFARX1 \key_mem_reg[7][89]  (.D(n4003), .SI(n8802), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[7][89] ), .QN(n8801));
   SDFFARX1 \key_mem_reg[8][89]  (.D(n4004), .SI(n8674), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[8][89] ), .QN(n8673));
   SDFFARX1 \key_mem_reg[9][89]  (.D(n4005), .SI(n8546), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[9][89] ), .QN(n8545));
   SDFFARX1 \key_mem_reg[10][89]  (.D(n4006), .SI(n8418), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[10][89] ), .QN(n8417));
   SDFFARX1 \key_mem_reg[11][89]  (.D(n4007), .SI(n8290), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[11][89] ), .QN(n8289));
   SDFFARX1 \key_mem_reg[12][89]  (.D(n4008), .SI(n8163), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[12][89] ), .QN(n8162));
   SDFFARX1 \key_mem_reg[13][89]  (.D(n4009), .SI(n8035), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[13][89] ), .QN(n8034));
   SDFFARX1 \key_mem_reg[14][89]  (.D(n4010), .SI(n7907), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(\key_mem[14][89] ), .QN(n7906));
   SDFFARX1 \prev_key1_reg_reg[88]  (.D(n5385), .SI(n7669), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7439), .Q(prev_key1_reg[88]), .QN(n3));
   SDFFARX1 \prev_key0_reg_reg[88]  (.D(n5512), .SI(n7780), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(prev_key0_reg[88]), .QN(n7779));
   SDFFARX1 \key_mem_reg[0][88]  (.D(n4011), .SI(n9698), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[0][88] ), .QN(n9697));
   SDFFARX1 \key_mem_reg[1][88]  (.D(n4012), .SI(n9570), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[1][88] ), .QN(n9569));
   SDFFARX1 \key_mem_reg[2][88]  (.D(n4013), .SI(n9442), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[2][88] ), .QN(n9441));
   SDFFARX1 \key_mem_reg[3][88]  (.D(n4014), .SI(n9314), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[3][88] ), .QN(n9313));
   SDFFARX1 \key_mem_reg[4][88]  (.D(n4015), .SI(n9187), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[4][88] ), .QN(n9186));
   SDFFARX1 \key_mem_reg[5][88]  (.D(n4016), .SI(n9059), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[5][88] ), .QN(n9058));
   SDFFARX1 \key_mem_reg[6][88]  (.D(n4017), .SI(n8931), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[6][88] ), .QN(n8930));
   SDFFARX1 \key_mem_reg[7][88]  (.D(n4018), .SI(n8803), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[7][88] ), .QN(n8802));
   SDFFARX1 \key_mem_reg[8][88]  (.D(n4019), .SI(n8675), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[8][88] ), .QN(n8674));
   SDFFARX1 \key_mem_reg[9][88]  (.D(n4020), .SI(n8547), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[9][88] ), .QN(n8546));
   SDFFARX1 \key_mem_reg[10][88]  (.D(n4021), .SI(n8419), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7438), .Q(\key_mem[10][88] ), .QN(n8418));
   SDFFARX1 \key_mem_reg[11][88]  (.D(n4022), .SI(n8291), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[11][88] ), .QN(n8290));
   SDFFARX1 \key_mem_reg[12][88]  (.D(n4023), .SI(n8164), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[12][88] ), .QN(n8163));
   SDFFARX1 \key_mem_reg[13][88]  (.D(n4024), .SI(n8036), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[13][88] ), .QN(n8035));
   SDFFARX1 \key_mem_reg[14][88]  (.D(n4025), .SI(n7908), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[14][88] ), .QN(n7907));
   SDFFARX1 \prev_key1_reg_reg[87]  (.D(n5386), .SI(n7670), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(prev_key1_reg[87]), .QN(n7669));
   SDFFARX1 \prev_key0_reg_reg[87]  (.D(n5513), .SI(n7781), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(prev_key0_reg[87]), .QN(n7780));
   SDFFARX1 \key_mem_reg[0][87]  (.D(n4026), .SI(n9699), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[0][87] ), .QN(n9698));
   SDFFARX1 \key_mem_reg[1][87]  (.D(n4027), .SI(n9571), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[1][87] ), .QN(n9570));
   SDFFARX1 \key_mem_reg[2][87]  (.D(n4028), .SI(n9443), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[2][87] ), .QN(n9442));
   SDFFARX1 \key_mem_reg[3][87]  (.D(n4029), .SI(n9315), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[3][87] ), .QN(n9314));
   SDFFARX1 \key_mem_reg[4][87]  (.D(n4030), .SI(n9188), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[4][87] ), .QN(n9187));
   SDFFARX1 \key_mem_reg[5][87]  (.D(n4031), .SI(n9060), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7437), .Q(\key_mem[5][87] ), .QN(n9059));
   SDFFARX1 \key_mem_reg[6][87]  (.D(n4032), .SI(n8932), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[6][87] ), .QN(n8931));
   SDFFARX1 \key_mem_reg[7][87]  (.D(n4033), .SI(n8804), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[7][87] ), .QN(n8803));
   SDFFARX1 \key_mem_reg[8][87]  (.D(n4034), .SI(n8676), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[8][87] ), .QN(n8675));
   SDFFARX1 \key_mem_reg[9][87]  (.D(n4035), .SI(n8548), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[9][87] ), .QN(n8547));
   SDFFARX1 \key_mem_reg[10][87]  (.D(n4036), .SI(n8420), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[10][87] ), .QN(n8419));
   SDFFARX1 \key_mem_reg[11][87]  (.D(n4037), .SI(n8292), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[11][87] ), .QN(n8291));
   SDFFARX1 \key_mem_reg[12][87]  (.D(n4038), .SI(n8165), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[12][87] ), .QN(n8164));
   SDFFARX1 \key_mem_reg[13][87]  (.D(n4039), .SI(n8037), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[13][87] ), .QN(n8036));
   SDFFARX1 \key_mem_reg[14][87]  (.D(n4040), .SI(n7909), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[14][87] ), .QN(n7908));
   SDFFARX1 \prev_key1_reg_reg[86]  (.D(n5387), .SI(n7671), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(prev_key1_reg[86]), .QN(n7670));
   SDFFARX1 \prev_key0_reg_reg[86]  (.D(n5514), .SI(n7782), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(prev_key0_reg[86]), .QN(n7781));
   SDFFARX1 \key_mem_reg[0][86]  (.D(n4041), .SI(n9700), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7436), .Q(\key_mem[0][86] ), .QN(n9699));
   SDFFARX1 \key_mem_reg[1][86]  (.D(n4042), .SI(n9572), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[1][86] ), .QN(n9571));
   SDFFARX1 \key_mem_reg[2][86]  (.D(n4043), .SI(n9444), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[2][86] ), .QN(n9443));
   SDFFARX1 \key_mem_reg[3][86]  (.D(n4044), .SI(n9316), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[3][86] ), .QN(n9315));
   SDFFARX1 \key_mem_reg[4][86]  (.D(n4045), .SI(n9189), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[4][86] ), .QN(n9188));
   SDFFARX1 \key_mem_reg[5][86]  (.D(n4046), .SI(n9061), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[5][86] ), .QN(n9060));
   SDFFARX1 \key_mem_reg[6][86]  (.D(n4047), .SI(n8933), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[6][86] ), .QN(n8932));
   SDFFARX1 \key_mem_reg[7][86]  (.D(n4048), .SI(n8805), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[7][86] ), .QN(n8804));
   SDFFARX1 \key_mem_reg[8][86]  (.D(n4049), .SI(n8677), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[8][86] ), .QN(n8676));
   SDFFARX1 \key_mem_reg[9][86]  (.D(n4050), .SI(n8549), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[9][86] ), .QN(n8548));
   SDFFARX1 \key_mem_reg[10][86]  (.D(n4051), .SI(n8421), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[10][86] ), .QN(n8420));
   SDFFARX1 \key_mem_reg[11][86]  (.D(n4052), .SI(n8293), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[11][86] ), .QN(n8292));
   SDFFARX1 \key_mem_reg[12][86]  (.D(n4053), .SI(n8166), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7435), .Q(\key_mem[12][86] ), .QN(n8165));
   SDFFARX1 \key_mem_reg[13][86]  (.D(n4054), .SI(n8038), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[13][86] ), .QN(n8037));
   SDFFARX1 \key_mem_reg[14][86]  (.D(n4055), .SI(n7910), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[14][86] ), .QN(n7909));
   SDFFARX1 \prev_key1_reg_reg[85]  (.D(n5388), .SI(n7672), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(prev_key1_reg[85]), .QN(n7671));
   SDFFARX1 \prev_key0_reg_reg[85]  (.D(n5515), .SI(n7783), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(prev_key0_reg[85]), .QN(n7782));
   SDFFARX1 \key_mem_reg[0][85]  (.D(n4056), .SI(n9701), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[0][85] ), .QN(n9700));
   SDFFARX1 \key_mem_reg[1][85]  (.D(n4057), .SI(n9573), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[1][85] ), .QN(n9572));
   SDFFARX1 \key_mem_reg[2][85]  (.D(n4058), .SI(n9445), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[2][85] ), .QN(n9444));
   SDFFARX1 \key_mem_reg[3][85]  (.D(n4059), .SI(n9317), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[3][85] ), .QN(n9316));
   SDFFARX1 \key_mem_reg[4][85]  (.D(n4060), .SI(n9190), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[4][85] ), .QN(n9189));
   SDFFARX1 \key_mem_reg[5][85]  (.D(n4061), .SI(n9062), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[5][85] ), .QN(n9061));
   SDFFARX1 \key_mem_reg[6][85]  (.D(n4062), .SI(n8934), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[6][85] ), .QN(n8933));
   SDFFARX1 \key_mem_reg[7][85]  (.D(n4063), .SI(n8806), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7434), .Q(\key_mem[7][85] ), .QN(n8805));
   SDFFARX1 \key_mem_reg[8][85]  (.D(n4064), .SI(n8678), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[8][85] ), .QN(n8677));
   SDFFARX1 \key_mem_reg[9][85]  (.D(n4065), .SI(n8550), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[9][85] ), .QN(n8549));
   SDFFARX1 \key_mem_reg[10][85]  (.D(n4066), .SI(n8422), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[10][85] ), .QN(n8421));
   SDFFARX1 \key_mem_reg[11][85]  (.D(n4067), .SI(n8294), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[11][85] ), .QN(n8293));
   SDFFARX1 \key_mem_reg[12][85]  (.D(n4068), .SI(n8167), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[12][85] ), .QN(n8166));
   SDFFARX1 \key_mem_reg[13][85]  (.D(n4069), .SI(n8039), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[13][85] ), .QN(n8038));
   SDFFARX1 \key_mem_reg[14][85]  (.D(n4070), .SI(n7911), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[14][85] ), .QN(n7910));
   SDFFARX1 \prev_key1_reg_reg[84]  (.D(n5389), .SI(n7673), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(prev_key1_reg[84]), .QN(n7672));
   SDFFARX1 \prev_key0_reg_reg[84]  (.D(n5516), .SI(n7784), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(prev_key0_reg[84]), .QN(n7783));
   SDFFARX1 \key_mem_reg[0][84]  (.D(n4071), .SI(n9702), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[0][84] ), .QN(n9701));
   SDFFARX1 \key_mem_reg[1][84]  (.D(n4072), .SI(n9574), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[1][84] ), .QN(n9573));
   SDFFARX1 \key_mem_reg[2][84]  (.D(n4073), .SI(n9446), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7433), .Q(\key_mem[2][84] ), .QN(n9445));
   SDFFARX1 \key_mem_reg[3][84]  (.D(n4074), .SI(n9318), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[3][84] ), .QN(n9317));
   SDFFARX1 \key_mem_reg[4][84]  (.D(n4075), .SI(n9191), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[4][84] ), .QN(n9190));
   SDFFARX1 \key_mem_reg[5][84]  (.D(n4076), .SI(n9063), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[5][84] ), .QN(n9062));
   SDFFARX1 \key_mem_reg[6][84]  (.D(n4077), .SI(n8935), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[6][84] ), .QN(n8934));
   SDFFARX1 \key_mem_reg[7][84]  (.D(n4078), .SI(n8807), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[7][84] ), .QN(n8806));
   SDFFARX1 \key_mem_reg[8][84]  (.D(n4079), .SI(n8679), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[8][84] ), .QN(n8678));
   SDFFARX1 \key_mem_reg[9][84]  (.D(n4080), .SI(n8551), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[9][84] ), .QN(n8550));
   SDFFARX1 \key_mem_reg[10][84]  (.D(n4081), .SI(n8423), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[10][84] ), .QN(n8422));
   SDFFARX1 \key_mem_reg[11][84]  (.D(n4082), .SI(n8295), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[11][84] ), .QN(n8294));
   SDFFARX1 \key_mem_reg[12][84]  (.D(n4083), .SI(n8168), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[12][84] ), .QN(n8167));
   SDFFARX1 \key_mem_reg[13][84]  (.D(n4084), .SI(n8040), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[13][84] ), .QN(n8039));
   SDFFARX1 \key_mem_reg[14][84]  (.D(n4085), .SI(n7912), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7432), .Q(\key_mem[14][84] ), .QN(n7911));
   SDFFARX1 \prev_key1_reg_reg[83]  (.D(n5390), .SI(n7674), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(prev_key1_reg[83]), .QN(n7673));
   SDFFARX1 \prev_key0_reg_reg[83]  (.D(n5517), .SI(n7785), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(prev_key0_reg[83]), .QN(n7784));
   SDFFARX1 \key_mem_reg[0][83]  (.D(n4086), .SI(n9703), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(\key_mem[0][83] ), .QN(n9702));
   SDFFARX1 \key_mem_reg[1][83]  (.D(n4087), .SI(n9575), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(\key_mem[1][83] ), .QN(n9574));
   SDFFARX1 \key_mem_reg[2][83]  (.D(n4088), .SI(n9447), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(\key_mem[2][83] ), .QN(n9446));
   SDFFARX1 \key_mem_reg[3][83]  (.D(n4089), .SI(n9319), .SE(test_se_buf_net1), .CLK(
          clk_buf_net1), .RSTB(n7431), .Q(\key_mem[3][83] ), .QN(n9318));
   SDFFARX1 \key_mem_reg[4][83]  (.D(n4090), .SI(n9192), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[4][83] ), .QN(n9191));
   SDFFARX1 \key_mem_reg[5][83]  (.D(n4091), .SI(n9064), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[5][83] ), .QN(n9063));
   SDFFARX1 \key_mem_reg[6][83]  (.D(n4092), .SI(n8936), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[6][83] ), .QN(n8935));
   SDFFARX1 \key_mem_reg[7][83]  (.D(n4093), .SI(n8808), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[7][83] ), .QN(n8807));
   SDFFARX1 \key_mem_reg[8][83]  (.D(n4094), .SI(n8680), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[8][83] ), .QN(n8679));
   SDFFARX1 \key_mem_reg[9][83]  (.D(n4095), .SI(n8552), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7431), .Q(\key_mem[9][83] ), .QN(n8551));
   SDFFARX1 \key_mem_reg[10][83]  (.D(n4096), .SI(n8424), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[10][83] ), .QN(n8423));
   SDFFARX1 \key_mem_reg[11][83]  (.D(n4097), .SI(n8296), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[11][83] ), .QN(n8295));
   SDFFARX1 \key_mem_reg[12][83]  (.D(n4098), .SI(n8169), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[12][83] ), .QN(n8168));
   SDFFARX1 \key_mem_reg[13][83]  (.D(n4099), .SI(n8041), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[13][83] ), .QN(n8040));
   SDFFARX1 \key_mem_reg[14][83]  (.D(n4100), .SI(n7913), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[14][83] ), .QN(n7912));
   SDFFARX1 \prev_key1_reg_reg[82]  (.D(n5391), .SI(n7675), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(prev_key1_reg[82]), .QN(n7674));
   SDFFARX1 \prev_key0_reg_reg[82]  (.D(n5518), .SI(n7786), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(prev_key0_reg[82]), .QN(n7785));
   SDFFARX1 \key_mem_reg[0][82]  (.D(n4101), .SI(n9704), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[0][82] ), .QN(n9703));
   SDFFARX1 \key_mem_reg[1][82]  (.D(n4102), .SI(n9576), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[1][82] ), .QN(n9575));
   SDFFARX1 \key_mem_reg[2][82]  (.D(n4103), .SI(n9448), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[2][82] ), .QN(n9447));
   SDFFARX1 \key_mem_reg[3][82]  (.D(n4104), .SI(n9320), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[3][82] ), .QN(n9319));
   SDFFARX1 \key_mem_reg[4][82]  (.D(n4105), .SI(n9193), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7430), .Q(\key_mem[4][82] ), .QN(n9192));
   SDFFARX1 \key_mem_reg[5][82]  (.D(n4106), .SI(n9065), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[5][82] ), .QN(n9064));
   SDFFARX1 \key_mem_reg[6][82]  (.D(n4107), .SI(n8937), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[6][82] ), .QN(n8936));
   SDFFARX1 \key_mem_reg[7][82]  (.D(n4108), .SI(n8809), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[7][82] ), .QN(n8808));
   SDFFARX1 \key_mem_reg[8][82]  (.D(n4109), .SI(n8681), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[8][82] ), .QN(n8680));
   SDFFARX1 \key_mem_reg[9][82]  (.D(n4110), .SI(n8553), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[9][82] ), .QN(n8552));
   SDFFARX1 \key_mem_reg[10][82]  (.D(n4111), .SI(n8425), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[10][82] ), .QN(n8424));
   SDFFARX1 \key_mem_reg[11][82]  (.D(n4112), .SI(n8297), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[11][82] ), .QN(n8296));
   SDFFARX1 \key_mem_reg[12][82]  (.D(n4113), .SI(n8170), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[12][82] ), .QN(n8169));
   SDFFARX1 \key_mem_reg[13][82]  (.D(n4114), .SI(n8042), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[13][82] ), .QN(n8041));
   SDFFARX1 \key_mem_reg[14][82]  (.D(n4115), .SI(n7914), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(\key_mem[14][82] ), .QN(n7913));
   SDFFARX1 \prev_key1_reg_reg[81]  (.D(n5392), .SI(n7676), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(prev_key1_reg[81]), .QN(n7675));
   SDFFARX1 \prev_key0_reg_reg[81]  (.D(n5519), .SI(n7787), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7429), .Q(prev_key0_reg[81]), .QN(n7786));
   SDFFARX1 \key_mem_reg[0][81]  (.D(n4116), .SI(n9705), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[0][81] ), .QN(n9704));
   SDFFARX1 \key_mem_reg[1][81]  (.D(n4117), .SI(n9577), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[1][81] ), .QN(n9576));
   SDFFARX1 \key_mem_reg[2][81]  (.D(n4118), .SI(n9449), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[2][81] ), .QN(n9448));
   SDFFARX1 \key_mem_reg[3][81]  (.D(n4119), .SI(n9321), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[3][81] ), .QN(n9320));
   SDFFARX1 \key_mem_reg[4][81]  (.D(n4120), .SI(n9194), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[4][81] ), .QN(n9193));
   SDFFARX1 \key_mem_reg[5][81]  (.D(n4121), .SI(n9066), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[5][81] ), .QN(n9065));
   SDFFARX1 \key_mem_reg[6][81]  (.D(n4122), .SI(n8938), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[6][81] ), .QN(n8937));
   SDFFARX1 \key_mem_reg[7][81]  (.D(n4123), .SI(n8810), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[7][81] ), .QN(n8809));
   SDFFARX1 \key_mem_reg[8][81]  (.D(n4124), .SI(n8682), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[8][81] ), .QN(n8681));
   SDFFARX1 \key_mem_reg[9][81]  (.D(n4125), .SI(n8554), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[9][81] ), .QN(n8553));
   SDFFARX1 \key_mem_reg[10][81]  (.D(n4126), .SI(n8426), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[10][81] ), .QN(n8425));
   SDFFARX1 \key_mem_reg[11][81]  (.D(n4127), .SI(n8298), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7428), .Q(\key_mem[11][81] ), .QN(n8297));
   SDFFARX1 \key_mem_reg[12][81]  (.D(n4128), .SI(n8171), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[12][81] ), .QN(n8170));
   SDFFARX1 \key_mem_reg[13][81]  (.D(n4129), .SI(n8043), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[13][81] ), .QN(n8042));
   SDFFARX1 \key_mem_reg[14][81]  (.D(n4130), .SI(n7915), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[14][81] ), .QN(n7914));
   SDFFARX1 \prev_key1_reg_reg[80]  (.D(n5393), .SI(n7677), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(prev_key1_reg[80]), .QN(n7676));
   SDFFARX1 \prev_key0_reg_reg[80]  (.D(n5520), .SI(n7788), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(prev_key0_reg[80]), .QN(n7787));
   SDFFARX1 \key_mem_reg[0][80]  (.D(n4131), .SI(n9706), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[0][80] ), .QN(n9705));
   SDFFARX1 \key_mem_reg[1][80]  (.D(n4132), .SI(n9578), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[1][80] ), .QN(n9577));
   SDFFARX1 \key_mem_reg[2][80]  (.D(n4133), .SI(n9450), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[2][80] ), .QN(n9449));
   SDFFARX1 \key_mem_reg[3][80]  (.D(n4134), .SI(n9322), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[3][80] ), .QN(n9321));
   SDFFARX1 \key_mem_reg[4][80]  (.D(n4135), .SI(n9195), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[4][80] ), .QN(n9194));
   SDFFARX1 \key_mem_reg[5][80]  (.D(n4136), .SI(n9067), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[5][80] ), .QN(n9066));
   SDFFARX1 \key_mem_reg[6][80]  (.D(n4137), .SI(n8939), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7427), .Q(\key_mem[6][80] ), .QN(n8938));
   SDFFARX1 \key_mem_reg[7][80]  (.D(n4138), .SI(n8811), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[7][80] ), .QN(n8810));
   SDFFARX1 \key_mem_reg[8][80]  (.D(n4139), .SI(n8683), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[8][80] ), .QN(n8682));
   SDFFARX1 \key_mem_reg[9][80]  (.D(n4140), .SI(n8555), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[9][80] ), .QN(n8554));
   SDFFARX1 \key_mem_reg[10][80]  (.D(n4141), .SI(n8427), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[10][80] ), .QN(n8426));
   SDFFARX1 \key_mem_reg[11][80]  (.D(n4142), .SI(n8299), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[11][80] ), .QN(n8298));
   SDFFARX1 \key_mem_reg[12][80]  (.D(n4143), .SI(n8172), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[12][80] ), .QN(n8171));
   SDFFARX1 \key_mem_reg[13][80]  (.D(n4144), .SI(n8044), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[13][80] ), .QN(n8043));
   SDFFARX1 \key_mem_reg[14][80]  (.D(n4145), .SI(n7916), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[14][80] ), .QN(n7915));
   SDFFARX1 \prev_key1_reg_reg[79]  (.D(n5394), .SI(n7678), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(prev_key1_reg[79]), .QN(n7677));
   SDFFARX1 \prev_key0_reg_reg[79]  (.D(n5521), .SI(n7789), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(prev_key0_reg[79]), .QN(n7788));
   SDFFARX1 \key_mem_reg[0][79]  (.D(n4146), .SI(n9707), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[0][79] ), .QN(n9706));
   SDFFARX1 \key_mem_reg[1][79]  (.D(n4147), .SI(n9579), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7426), .Q(\key_mem[1][79] ), .QN(n9578));
   SDFFARX1 \key_mem_reg[2][79]  (.D(n4148), .SI(n9451), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[2][79] ), .QN(n9450));
   SDFFARX1 \key_mem_reg[3][79]  (.D(n4149), .SI(n9323), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[3][79] ), .QN(n9322));
   SDFFARX1 \key_mem_reg[4][79]  (.D(n4150), .SI(n9196), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[4][79] ), .QN(n9195));
   SDFFARX1 \key_mem_reg[5][79]  (.D(n4151), .SI(n9068), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[5][79] ), .QN(n9067));
   SDFFARX1 \key_mem_reg[6][79]  (.D(n4152), .SI(n8940), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[6][79] ), .QN(n8939));
   SDFFARX1 \key_mem_reg[7][79]  (.D(n4153), .SI(n8812), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[7][79] ), .QN(n8811));
   SDFFARX1 \key_mem_reg[8][79]  (.D(n4154), .SI(n8684), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[8][79] ), .QN(n8683));
   SDFFARX1 \key_mem_reg[9][79]  (.D(n4155), .SI(n8556), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[9][79] ), .QN(n8555));
   SDFFARX1 \key_mem_reg[10][79]  (.D(n4156), .SI(n8428), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[10][79] ), .QN(n8427));
   SDFFARX1 \key_mem_reg[11][79]  (.D(n4157), .SI(n8300), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[11][79] ), .QN(n8299));
   SDFFARX1 \key_mem_reg[12][79]  (.D(n4158), .SI(n8173), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[12][79] ), .QN(n8172));
   SDFFARX1 \key_mem_reg[13][79]  (.D(n4159), .SI(n8045), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7425), .Q(\key_mem[13][79] ), .QN(n8044));
   SDFFARX1 \key_mem_reg[14][79]  (.D(n4160), .SI(n7917), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[14][79] ), .QN(n7916));
   SDFFARX1 \prev_key1_reg_reg[78]  (.D(n5395), .SI(n7679), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(prev_key1_reg[78]), .QN(n7678));
   SDFFARX1 \prev_key0_reg_reg[78]  (.D(n5522), .SI(n7790), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(prev_key0_reg[78]), .QN(n7789));
   SDFFARX1 \key_mem_reg[0][78]  (.D(n4161), .SI(n9708), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[0][78] ), .QN(n9707));
   SDFFARX1 \key_mem_reg[1][78]  (.D(n4162), .SI(n9580), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[1][78] ), .QN(n9579));
   SDFFARX1 \key_mem_reg[2][78]  (.D(n4163), .SI(n9452), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[2][78] ), .QN(n9451));
   SDFFARX1 \key_mem_reg[3][78]  (.D(n4164), .SI(n9324), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[3][78] ), .QN(n9323));
   SDFFARX1 \key_mem_reg[4][78]  (.D(n4165), .SI(test_si2), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[4][78] ), .QN(n9196));
   SDFFARX1 \key_mem_reg[5][78]  (.D(n4166), .SI(n9069), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[5][78] ), .QN(n9068));
   SDFFARX1 \key_mem_reg[6][78]  (.D(n4167), .SI(n8941), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[6][78] ), .QN(n8940));
   SDFFARX1 \key_mem_reg[7][78]  (.D(n4168), .SI(n8813), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[7][78] ), .QN(n8812));
   SDFFARX1 \key_mem_reg[8][78]  (.D(n4169), .SI(n8685), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7424), .Q(\key_mem[8][78] ), .QN(n8684));
   SDFFARX1 \key_mem_reg[9][78]  (.D(n4170), .SI(n8557), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[9][78] ), .QN(n8556));
   SDFFARX1 \key_mem_reg[10][78]  (.D(n4171), .SI(n8429), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[10][78] ), .QN(n8428));
   SDFFARX1 \key_mem_reg[11][78]  (.D(n4172), .SI(n8301), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[11][78] ), .QN(n8300));
   SDFFARX1 \key_mem_reg[12][78]  (.D(n4173), .SI(n8174), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[12][78] ), .QN(n8173));
   SDFFARX1 \key_mem_reg[13][78]  (.D(n4174), .SI(n8046), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[13][78] ), .QN(n8045));
   SDFFARX1 \key_mem_reg[14][78]  (.D(n4175), .SI(n7918), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[14][78] ), .QN(n7917));
   SDFFARX1 \prev_key1_reg_reg[77]  (.D(n5396), .SI(n7680), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(prev_key1_reg[77]), .QN(n7679));
   SDFFARX1 \prev_key0_reg_reg[77]  (.D(n5523), .SI(n7791), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(prev_key0_reg[77]), .QN(n7790));
   SDFFARX1 \key_mem_reg[0][77]  (.D(n4176), .SI(n9709), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[0][77] ), .QN(n9708));
   SDFFARX1 \key_mem_reg[1][77]  (.D(n4177), .SI(n9581), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[1][77] ), .QN(n9580));
   SDFFARX1 \key_mem_reg[2][77]  (.D(n4178), .SI(n9453), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[2][77] ), .QN(n9452));
   SDFFARX1 \key_mem_reg[3][77]  (.D(n4179), .SI(n9325), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7423), .Q(\key_mem[3][77] ), .QN(n9324));
   SDFFARX1 \key_mem_reg[4][77]  (.D(n4180), .SI(n9197), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[4][77] ));
   SDFFARX1 \key_mem_reg[5][77]  (.D(n4181), .SI(n9070), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[5][77] ), .QN(n9069));
   SDFFARX1 \key_mem_reg[6][77]  (.D(n4182), .SI(n8942), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[6][77] ), .QN(n8941));
   SDFFARX1 \key_mem_reg[7][77]  (.D(n4183), .SI(n8814), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[7][77] ), .QN(n8813));
   SDFFARX1 \key_mem_reg[8][77]  (.D(n4184), .SI(n8686), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[8][77] ), .QN(n8685));
   SDFFARX1 \key_mem_reg[9][77]  (.D(n4185), .SI(n8558), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[9][77] ), .QN(n8557));
   SDFFARX1 \key_mem_reg[10][77]  (.D(n4186), .SI(n8430), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[10][77] ), .QN(n8429));
   SDFFARX1 \key_mem_reg[11][77]  (.D(n4187), .SI(n8302), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[11][77] ), .QN(n8301));
   SDFFARX1 \key_mem_reg[12][77]  (.D(n4188), .SI(n8175), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[12][77] ), .QN(n8174));
   SDFFARX1 \key_mem_reg[13][77]  (.D(n4189), .SI(n8047), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[13][77] ), .QN(n8046));
   SDFFARX1 \key_mem_reg[14][77]  (.D(n4190), .SI(n7919), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(\key_mem[14][77] ), .QN(n7918));
   SDFFARX1 \prev_key1_reg_reg[76]  (.D(n5397), .SI(n7681), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7422), .Q(prev_key1_reg[76]), .QN(n7680));
   SDFFARX1 \prev_key0_reg_reg[76]  (.D(n5524), .SI(n7792), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(prev_key0_reg[76]), .QN(n7791));
   SDFFARX1 \key_mem_reg[0][76]  (.D(n4191), .SI(n9710), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[0][76] ), .QN(n9709));
   SDFFARX1 \key_mem_reg[1][76]  (.D(n4192), .SI(n9582), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[1][76] ), .QN(n9581));
   SDFFARX1 \key_mem_reg[2][76]  (.D(n4193), .SI(n9454), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[2][76] ), .QN(n9453));
   SDFFARX1 \key_mem_reg[3][76]  (.D(n4194), .SI(n9326), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[3][76] ), .QN(n9325));
   SDFFARX1 \key_mem_reg[4][76]  (.D(n4195), .SI(n9198), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[4][76] ), .QN(n9197));
   SDFFARX1 \key_mem_reg[5][76]  (.D(n4196), .SI(n9071), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[5][76] ), .QN(n9070));
   SDFFARX1 \key_mem_reg[6][76]  (.D(n4197), .SI(n8943), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[6][76] ), .QN(n8942));
   SDFFARX1 \key_mem_reg[7][76]  (.D(n4198), .SI(n8815), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[7][76] ), .QN(n8814));
   SDFFARX1 \key_mem_reg[8][76]  (.D(n4199), .SI(n8687), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[8][76] ), .QN(n8686));
   SDFFARX1 \key_mem_reg[9][76]  (.D(n4200), .SI(n8559), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[9][76] ), .QN(n8558));
   SDFFARX1 \key_mem_reg[10][76]  (.D(n4201), .SI(n8431), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7421), .Q(\key_mem[10][76] ), .QN(n8430));
   SDFFARX1 \key_mem_reg[11][76]  (.D(n4202), .SI(n8303), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[11][76] ), .QN(n8302));
   SDFFARX1 \key_mem_reg[12][76]  (.D(n4203), .SI(n8176), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[12][76] ), .QN(n8175));
   SDFFARX1 \key_mem_reg[13][76]  (.D(n4204), .SI(n8048), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[13][76] ), .QN(n8047));
   SDFFARX1 \key_mem_reg[14][76]  (.D(n4205), .SI(n7920), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[14][76] ), .QN(n7919));
   SDFFARX1 \prev_key1_reg_reg[75]  (.D(n5398), .SI(n7682), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(prev_key1_reg[75]), .QN(n7681));
   SDFFARX1 \prev_key0_reg_reg[75]  (.D(n5525), .SI(n7793), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(prev_key0_reg[75]), .QN(n7792));
   SDFFARX1 \key_mem_reg[0][75]  (.D(n4206), .SI(n9711), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[0][75] ), .QN(n9710));
   SDFFARX1 \key_mem_reg[1][75]  (.D(n4207), .SI(n9583), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[1][75] ), .QN(n9582));
   SDFFARX1 \key_mem_reg[2][75]  (.D(n4208), .SI(n9455), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[2][75] ), .QN(n9454));
   SDFFARX1 \key_mem_reg[3][75]  (.D(n4209), .SI(n9327), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[3][75] ), .QN(n9326));
   SDFFARX1 \key_mem_reg[4][75]  (.D(n4210), .SI(n9199), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[4][75] ), .QN(n9198));
   SDFFARX1 \key_mem_reg[5][75]  (.D(n4211), .SI(n9072), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7420), .Q(\key_mem[5][75] ), .QN(n9071));
   SDFFARX1 \key_mem_reg[6][75]  (.D(n4212), .SI(n8944), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[6][75] ), .QN(n8943));
   SDFFARX1 \key_mem_reg[7][75]  (.D(n4213), .SI(n8816), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[7][75] ), .QN(n8815));
   SDFFARX1 \key_mem_reg[8][75]  (.D(n4214), .SI(n8688), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[8][75] ), .QN(n8687));
   SDFFARX1 \key_mem_reg[9][75]  (.D(n4215), .SI(n8560), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[9][75] ), .QN(n8559));
   SDFFARX1 \key_mem_reg[10][75]  (.D(n4216), .SI(n8432), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[10][75] ), .QN(n8431));
   SDFFARX1 \key_mem_reg[11][75]  (.D(n4217), .SI(n8304), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[11][75] ), .QN(n8303));
   SDFFARX1 \key_mem_reg[12][75]  (.D(n4218), .SI(n8177), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[12][75] ), .QN(n8176));
   SDFFARX1 \key_mem_reg[13][75]  (.D(n4219), .SI(n8049), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[13][75] ), .QN(n8048));
   SDFFARX1 \key_mem_reg[14][75]  (.D(n4220), .SI(n7921), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[14][75] ), .QN(n7920));
   SDFFARX1 \prev_key1_reg_reg[74]  (.D(n5399), .SI(n7683), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(prev_key1_reg[74]), .QN(n7682));
   SDFFARX1 \prev_key0_reg_reg[74]  (.D(n5526), .SI(n7794), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(prev_key0_reg[74]), .QN(n7793));
   SDFFARX1 \key_mem_reg[0][74]  (.D(n4221), .SI(n9712), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7419), .Q(\key_mem[0][74] ), .QN(n9711));
   SDFFARX1 \key_mem_reg[1][74]  (.D(n4222), .SI(n9584), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[1][74] ), .QN(n9583));
   SDFFARX1 \key_mem_reg[2][74]  (.D(n4223), .SI(n9456), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[2][74] ), .QN(n9455));
   SDFFARX1 \key_mem_reg[3][74]  (.D(n4224), .SI(n9328), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[3][74] ), .QN(n9327));
   SDFFARX1 \key_mem_reg[4][74]  (.D(n4225), .SI(n9200), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[4][74] ), .QN(n9199));
   SDFFARX1 \key_mem_reg[5][74]  (.D(n4226), .SI(n9073), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[5][74] ), .QN(n9072));
   SDFFARX1 \key_mem_reg[6][74]  (.D(n4227), .SI(n8945), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[6][74] ), .QN(n8944));
   SDFFARX1 \key_mem_reg[7][74]  (.D(n4228), .SI(n8817), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[7][74] ), .QN(n8816));
   SDFFARX1 \key_mem_reg[8][74]  (.D(n4229), .SI(n8689), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[8][74] ), .QN(n8688));
   SDFFARX1 \key_mem_reg[9][74]  (.D(n4230), .SI(n8561), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[9][74] ), .QN(n8560));
   SDFFARX1 \key_mem_reg[10][74]  (.D(n4231), .SI(n8433), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[10][74] ), .QN(n8432));
   SDFFARX1 \key_mem_reg[11][74]  (.D(n4232), .SI(n8305), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[11][74] ), .QN(n8304));
   SDFFARX1 \key_mem_reg[12][74]  (.D(n4233), .SI(n8178), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7418), .Q(\key_mem[12][74] ), .QN(n8177));
   SDFFARX1 \key_mem_reg[13][74]  (.D(n4234), .SI(n8050), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[13][74] ), .QN(n8049));
   SDFFARX1 \key_mem_reg[14][74]  (.D(n4235), .SI(n7922), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[14][74] ), .QN(n7921));
   SDFFARX1 \prev_key1_reg_reg[73]  (.D(n5400), .SI(n7684), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(prev_key1_reg[73]), .QN(n7683));
   SDFFARX1 \prev_key0_reg_reg[73]  (.D(n5527), .SI(n7795), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(prev_key0_reg[73]), .QN(n7794));
   SDFFARX1 \key_mem_reg[0][73]  (.D(n4236), .SI(n9713), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[0][73] ), .QN(n9712));
   SDFFARX1 \key_mem_reg[1][73]  (.D(n4237), .SI(n9585), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[1][73] ), .QN(n9584));
   SDFFARX1 \key_mem_reg[2][73]  (.D(n4238), .SI(n9457), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[2][73] ), .QN(n9456));
   SDFFARX1 \key_mem_reg[3][73]  (.D(n4239), .SI(n9329), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[3][73] ), .QN(n9328));
   SDFFARX1 \key_mem_reg[4][73]  (.D(n4240), .SI(n9201), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[4][73] ), .QN(n9200));
   SDFFARX1 \key_mem_reg[5][73]  (.D(n4241), .SI(n9074), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[5][73] ), .QN(n9073));
   SDFFARX1 \key_mem_reg[6][73]  (.D(n4242), .SI(n8946), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[6][73] ), .QN(n8945));
   SDFFARX1 \key_mem_reg[7][73]  (.D(n4243), .SI(n8818), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7417), .Q(\key_mem[7][73] ), .QN(n8817));
   SDFFARX1 \key_mem_reg[8][73]  (.D(n4244), .SI(n8690), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[8][73] ), .QN(n8689));
   SDFFARX1 \key_mem_reg[9][73]  (.D(n4245), .SI(n8562), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[9][73] ), .QN(n8561));
   SDFFARX1 \key_mem_reg[10][73]  (.D(n4246), .SI(n8434), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[10][73] ), .QN(n8433));
   SDFFARX1 \key_mem_reg[11][73]  (.D(n4247), .SI(n8306), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[11][73] ), .QN(n8305));
   SDFFARX1 \key_mem_reg[12][73]  (.D(n4248), .SI(n8179), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[12][73] ), .QN(n8178));
   SDFFARX1 \key_mem_reg[13][73]  (.D(n4249), .SI(n8051), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[13][73] ), .QN(n8050));
   SDFFARX1 \key_mem_reg[14][73]  (.D(n4250), .SI(n7923), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[14][73] ), .QN(n7922));
   SDFFARX1 \prev_key1_reg_reg[72]  (.D(n5401), .SI(n7685), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(prev_key1_reg[72]), .QN(n7684));
   SDFFARX1 \prev_key0_reg_reg[72]  (.D(n5528), .SI(n7796), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(prev_key0_reg[72]), .QN(n7795));
   SDFFARX1 \key_mem_reg[0][72]  (.D(n4251), .SI(n9714), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[0][72] ), .QN(n9713));
   SDFFARX1 \key_mem_reg[1][72]  (.D(n4252), .SI(n9586), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[1][72] ), .QN(n9585));
   SDFFARX1 \key_mem_reg[2][72]  (.D(n4253), .SI(n9458), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7416), .Q(\key_mem[2][72] ), .QN(n9457));
   SDFFARX1 \key_mem_reg[3][72]  (.D(n4254), .SI(n9330), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[3][72] ), .QN(n9329));
   SDFFARX1 \key_mem_reg[4][72]  (.D(n4255), .SI(n9202), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[4][72] ), .QN(n9201));
   SDFFARX1 \key_mem_reg[5][72]  (.D(n4256), .SI(n9075), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[5][72] ), .QN(n9074));
   SDFFARX1 \key_mem_reg[6][72]  (.D(n4257), .SI(n8947), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[6][72] ), .QN(n8946));
   SDFFARX1 \key_mem_reg[7][72]  (.D(n4258), .SI(n8819), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[7][72] ), .QN(n8818));
   SDFFARX1 \key_mem_reg[8][72]  (.D(n4259), .SI(n8691), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[8][72] ), .QN(n8690));
   SDFFARX1 \key_mem_reg[9][72]  (.D(n4260), .SI(n8563), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[9][72] ), .QN(n8562));
   SDFFARX1 \key_mem_reg[10][72]  (.D(n4261), .SI(n8435), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[10][72] ), .QN(n8434));
   SDFFARX1 \key_mem_reg[11][72]  (.D(n4262), .SI(n8307), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[11][72] ), .QN(n8306));
   SDFFARX1 \key_mem_reg[12][72]  (.D(n4263), .SI(n8180), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[12][72] ), .QN(n8179));
   SDFFARX1 \key_mem_reg[13][72]  (.D(n4264), .SI(n8052), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[13][72] ), .QN(n8051));
   SDFFARX1 \key_mem_reg[14][72]  (.D(n4265), .SI(n7924), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7415), .Q(\key_mem[14][72] ), .QN(n7923));
   SDFFARX1 \prev_key1_reg_reg[71]  (.D(n5402), .SI(n7686), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(prev_key1_reg[71]), .QN(n7685));
   SDFFARX1 \prev_key0_reg_reg[71]  (.D(n5529), .SI(n7797), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(prev_key0_reg[71]), .QN(n7796));
   SDFFARX1 \key_mem_reg[0][71]  (.D(n4266), .SI(n9715), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[0][71] ), .QN(n9714));
   SDFFARX1 \key_mem_reg[1][71]  (.D(n4267), .SI(n9587), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[1][71] ), .QN(n9586));
   SDFFARX1 \key_mem_reg[2][71]  (.D(n4268), .SI(n9459), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[2][71] ), .QN(n9458));
   SDFFARX1 \key_mem_reg[3][71]  (.D(n4269), .SI(n9331), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[3][71] ), .QN(n9330));
   SDFFARX1 \key_mem_reg[4][71]  (.D(n4270), .SI(n9203), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[4][71] ), .QN(n9202));
   SDFFARX1 \key_mem_reg[5][71]  (.D(n4271), .SI(n9076), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[5][71] ), .QN(n9075));
   SDFFARX1 \key_mem_reg[6][71]  (.D(n4272), .SI(n8948), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[6][71] ), .QN(n8947));
   SDFFARX1 \key_mem_reg[7][71]  (.D(n4273), .SI(n8820), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[7][71] ), .QN(n8819));
   SDFFARX1 \key_mem_reg[8][71]  (.D(n4274), .SI(n8692), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[8][71] ), .QN(n8691));
   SDFFARX1 \key_mem_reg[9][71]  (.D(n4275), .SI(n8564), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7414), .Q(\key_mem[9][71] ), .QN(n8563));
   SDFFARX1 \key_mem_reg[10][71]  (.D(n4276), .SI(n8436), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[10][71] ), .QN(n8435));
   SDFFARX1 \key_mem_reg[11][71]  (.D(n4277), .SI(n8308), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[11][71] ), .QN(n8307));
   SDFFARX1 \key_mem_reg[12][71]  (.D(n4278), .SI(n8181), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[12][71] ), .QN(n8180));
   SDFFARX1 \key_mem_reg[13][71]  (.D(n4279), .SI(n8053), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[13][71] ), .QN(n8052));
   SDFFARX1 \key_mem_reg[14][71]  (.D(n4280), .SI(n7925), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[14][71] ), .QN(n7924));
   SDFFARX1 \prev_key1_reg_reg[70]  (.D(n5403), .SI(n7687), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(prev_key1_reg[70]), .QN(n7686));
   SDFFARX1 \prev_key0_reg_reg[70]  (.D(n5530), .SI(n7798), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(prev_key0_reg[70]), .QN(n7797));
   SDFFARX1 \key_mem_reg[0][70]  (.D(n4281), .SI(n9716), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[0][70] ), .QN(n9715));
   SDFFARX1 \key_mem_reg[1][70]  (.D(n4282), .SI(n9588), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[1][70] ), .QN(n9587));
   SDFFARX1 \key_mem_reg[2][70]  (.D(n4283), .SI(n9460), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[2][70] ), .QN(n9459));
   SDFFARX1 \key_mem_reg[3][70]  (.D(n4284), .SI(n9332), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[3][70] ), .QN(n9331));
   SDFFARX1 \key_mem_reg[4][70]  (.D(n4285), .SI(n9204), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7413), .Q(\key_mem[4][70] ), .QN(n9203));
   SDFFARX1 \key_mem_reg[5][70]  (.D(n4286), .SI(n9077), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[5][70] ), .QN(n9076));
   SDFFARX1 \key_mem_reg[6][70]  (.D(n4287), .SI(n8949), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[6][70] ), .QN(n8948));
   SDFFARX1 \key_mem_reg[7][70]  (.D(n4288), .SI(n8821), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[7][70] ), .QN(n8820));
   SDFFARX1 \key_mem_reg[8][70]  (.D(n4289), .SI(n8693), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[8][70] ), .QN(n8692));
   SDFFARX1 \key_mem_reg[9][70]  (.D(n4290), .SI(n8565), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[9][70] ), .QN(n8564));
   SDFFARX1 \key_mem_reg[10][70]  (.D(n4291), .SI(n8437), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[10][70] ), .QN(n8436));
   SDFFARX1 \key_mem_reg[11][70]  (.D(n4292), .SI(n8309), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[11][70] ), .QN(n8308));
   SDFFARX1 \key_mem_reg[12][70]  (.D(n4293), .SI(n8182), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[12][70] ), .QN(n8181));
   SDFFARX1 \key_mem_reg[13][70]  (.D(n4294), .SI(n8054), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[13][70] ), .QN(n8053));
   SDFFARX1 \key_mem_reg[14][70]  (.D(n4295), .SI(n7926), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(\key_mem[14][70] ), .QN(n7925));
   SDFFARX1 \prev_key1_reg_reg[69]  (.D(n5404), .SI(n7688), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(prev_key1_reg[69]), .QN(n7687));
   SDFFARX1 \prev_key0_reg_reg[69]  (.D(n5531), .SI(n7799), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7412), .Q(prev_key0_reg[69]), .QN(n7798));
   SDFFARX1 \key_mem_reg[0][69]  (.D(n4296), .SI(n9717), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[0][69] ), .QN(n9716));
   SDFFARX1 \key_mem_reg[1][69]  (.D(n4297), .SI(n9589), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[1][69] ), .QN(n9588));
   SDFFARX1 \key_mem_reg[2][69]  (.D(n4298), .SI(n9461), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[2][69] ), .QN(n9460));
   SDFFARX1 \key_mem_reg[3][69]  (.D(n4299), .SI(n9333), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[3][69] ), .QN(n9332));
   SDFFARX1 \key_mem_reg[4][69]  (.D(n4300), .SI(n9205), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[4][69] ), .QN(n9204));
   SDFFARX1 \key_mem_reg[5][69]  (.D(n4301), .SI(n9078), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[5][69] ), .QN(n9077));
   SDFFARX1 \key_mem_reg[6][69]  (.D(n4302), .SI(n8950), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[6][69] ), .QN(n8949));
   SDFFARX1 \key_mem_reg[7][69]  (.D(n4303), .SI(n8822), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[7][69] ), .QN(n8821));
   SDFFARX1 \key_mem_reg[8][69]  (.D(n4304), .SI(n8694), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[8][69] ), .QN(n8693));
   SDFFARX1 \key_mem_reg[9][69]  (.D(n4305), .SI(n8566), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[9][69] ), .QN(n8565));
   SDFFARX1 \key_mem_reg[10][69]  (.D(n4306), .SI(n8438), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[10][69] ), .QN(n8437));
   SDFFARX1 \key_mem_reg[11][69]  (.D(n4307), .SI(n8310), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7411), .Q(\key_mem[11][69] ), .QN(n8309));
   SDFFARX1 \key_mem_reg[12][69]  (.D(n4308), .SI(n8183), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[12][69] ), .QN(n8182));
   SDFFARX1 \key_mem_reg[13][69]  (.D(n4309), .SI(n8055), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[13][69] ), .QN(n8054));
   SDFFARX1 \key_mem_reg[14][69]  (.D(n4310), .SI(n7927), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[14][69] ), .QN(n7926));
   SDFFARX1 \prev_key1_reg_reg[68]  (.D(n5405), .SI(n7689), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(prev_key1_reg[68]), .QN(n7688));
   SDFFARX1 \prev_key0_reg_reg[68]  (.D(n5532), .SI(n7800), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(prev_key0_reg[68]), .QN(n7799));
   SDFFARX1 \key_mem_reg[0][68]  (.D(n4311), .SI(n9718), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[0][68] ), .QN(n9717));
   SDFFARX1 \key_mem_reg[1][68]  (.D(n4312), .SI(n9590), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[1][68] ), .QN(n9589));
   SDFFARX1 \key_mem_reg[2][68]  (.D(n4313), .SI(n9462), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[2][68] ), .QN(n9461));
   SDFFARX1 \key_mem_reg[3][68]  (.D(n4314), .SI(n9334), .SE(test_se_buf_net2), .CLK(
          clk_buf_net2), .RSTB(n7410), .Q(\key_mem[3][68] ), .QN(n9333));
   SDFFARX1 \key_mem_reg[4][68]  (.D(n4315), .SI(n9206), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7410), .Q(\key_mem[4][68] ), .QN(n9205));
   SDFFARX1 \key_mem_reg[5][68]  (.D(n4316), .SI(n9079), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7410), .Q(\key_mem[5][68] ), .QN(n9078));
   SDFFARX1 \key_mem_reg[6][68]  (.D(n4317), .SI(n8951), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7410), .Q(\key_mem[6][68] ), .QN(n8950));
   SDFFARX1 \key_mem_reg[7][68]  (.D(n4318), .SI(n8823), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[7][68] ), .QN(n8822));
   SDFFARX1 \key_mem_reg[8][68]  (.D(n4319), .SI(n8695), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[8][68] ), .QN(n8694));
   SDFFARX1 \key_mem_reg[9][68]  (.D(n4320), .SI(n8567), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[9][68] ), .QN(n8566));
   SDFFARX1 \key_mem_reg[10][68]  (.D(n4321), .SI(n8439), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[10][68] ), .QN(n8438));
   SDFFARX1 \key_mem_reg[11][68]  (.D(n4322), .SI(n8311), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[11][68] ), .QN(n8310));
   SDFFARX1 \key_mem_reg[12][68]  (.D(n4323), .SI(n8184), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[12][68] ), .QN(n8183));
   SDFFARX1 \key_mem_reg[13][68]  (.D(n4324), .SI(n8056), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[13][68] ), .QN(n8055));
   SDFFARX1 \key_mem_reg[14][68]  (.D(n4325), .SI(n7928), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[14][68] ), .QN(n7927));
   SDFFARX1 \prev_key1_reg_reg[67]  (.D(n5406), .SI(n7690), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(prev_key1_reg[67]), .QN(n7689));
   SDFFARX1 \prev_key0_reg_reg[67]  (.D(n5533), .SI(n7801), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(prev_key0_reg[67]), .QN(n7800));
   SDFFARX1 \key_mem_reg[0][67]  (.D(n4326), .SI(n9719), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[0][67] ), .QN(n9718));
   SDFFARX1 \key_mem_reg[1][67]  (.D(n4327), .SI(n9591), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7409), .Q(\key_mem[1][67] ), .QN(n9590));
   SDFFARX1 \key_mem_reg[2][67]  (.D(n4328), .SI(n9463), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[2][67] ), .QN(n9462));
   SDFFARX1 \key_mem_reg[3][67]  (.D(n4329), .SI(n9335), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[3][67] ), .QN(n9334));
   SDFFARX1 \key_mem_reg[4][67]  (.D(n4330), .SI(n9207), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[4][67] ), .QN(n9206));
   SDFFARX1 \key_mem_reg[5][67]  (.D(n4331), .SI(n9080), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[5][67] ), .QN(n9079));
   SDFFARX1 \key_mem_reg[6][67]  (.D(n4332), .SI(n8952), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[6][67] ), .QN(n8951));
   SDFFARX1 \key_mem_reg[7][67]  (.D(n4333), .SI(n8824), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[7][67] ), .QN(n8823));
   SDFFARX1 \key_mem_reg[8][67]  (.D(n4334), .SI(n8696), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[8][67] ), .QN(n8695));
   SDFFARX1 \key_mem_reg[9][67]  (.D(n4335), .SI(n8568), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[9][67] ), .QN(n8567));
   SDFFARX1 \key_mem_reg[10][67]  (.D(n4336), .SI(n8440), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[10][67] ), .QN(n8439));
   SDFFARX1 \key_mem_reg[11][67]  (.D(n4337), .SI(n8312), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[11][67] ), .QN(n8311));
   SDFFARX1 \key_mem_reg[12][67]  (.D(n4338), .SI(n8185), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[12][67] ), .QN(n8184));
   SDFFARX1 \key_mem_reg[13][67]  (.D(n4339), .SI(n8057), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7408), .Q(\key_mem[13][67] ), .QN(n8056));
   SDFFARX1 \key_mem_reg[14][67]  (.D(n4340), .SI(n7929), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[14][67] ), .QN(n7928));
   SDFFARX1 \prev_key1_reg_reg[66]  (.D(n5407), .SI(n7691), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(prev_key1_reg[66]), .QN(n7690));
   SDFFARX1 \prev_key0_reg_reg[66]  (.D(n5534), .SI(n7802), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(prev_key0_reg[66]), .QN(n7801));
   SDFFARX1 \key_mem_reg[0][66]  (.D(n4341), .SI(n9720), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[0][66] ), .QN(n9719));
   SDFFARX1 \key_mem_reg[1][66]  (.D(n4342), .SI(n9592), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[1][66] ), .QN(n9591));
   SDFFARX1 \key_mem_reg[2][66]  (.D(n4343), .SI(n9464), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[2][66] ), .QN(n9463));
   SDFFARX1 \key_mem_reg[3][66]  (.D(n4344), .SI(n9336), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[3][66] ), .QN(n9335));
   SDFFARX1 \key_mem_reg[4][66]  (.D(n4345), .SI(n9208), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[4][66] ), .QN(n9207));
   SDFFARX1 \key_mem_reg[5][66]  (.D(n4346), .SI(n9081), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[5][66] ), .QN(n9080));
   SDFFARX1 \key_mem_reg[6][66]  (.D(n4347), .SI(n8953), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[6][66] ), .QN(n8952));
   SDFFARX1 \key_mem_reg[7][66]  (.D(n4348), .SI(n8825), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[7][66] ), .QN(n8824));
   SDFFARX1 \key_mem_reg[8][66]  (.D(n4349), .SI(n8697), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7407), .Q(\key_mem[8][66] ), .QN(n8696));
   SDFFARX1 \key_mem_reg[9][66]  (.D(n4350), .SI(n8569), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[9][66] ), .QN(n8568));
   SDFFARX1 \key_mem_reg[10][66]  (.D(n4351), .SI(n8441), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[10][66] ), .QN(n8440));
   SDFFARX1 \key_mem_reg[11][66]  (.D(n4352), .SI(n8313), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[11][66] ), .QN(n8312));
   SDFFARX1 \key_mem_reg[12][66]  (.D(n4353), .SI(n8186), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[12][66] ), .QN(n8185));
   SDFFARX1 \key_mem_reg[13][66]  (.D(n4354), .SI(n8058), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[13][66] ), .QN(n8057));
   SDFFARX1 \key_mem_reg[14][66]  (.D(n4355), .SI(n7930), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[14][66] ), .QN(n7929));
   SDFFARX1 \prev_key1_reg_reg[65]  (.D(n5408), .SI(n7692), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(prev_key1_reg[65]), .QN(n7691));
   SDFFARX1 \prev_key0_reg_reg[65]  (.D(n5535), .SI(n7803), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(prev_key0_reg[65]), .QN(n7802));
   SDFFARX1 \key_mem_reg[0][65]  (.D(n4356), .SI(n9721), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[0][65] ), .QN(n9720));
   SDFFARX1 \key_mem_reg[1][65]  (.D(n4357), .SI(n9593), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[1][65] ), .QN(n9592));
   SDFFARX1 \key_mem_reg[2][65]  (.D(n4358), .SI(n9465), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[2][65] ), .QN(n9464));
   SDFFARX1 \key_mem_reg[3][65]  (.D(n4359), .SI(n9337), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7406), .Q(\key_mem[3][65] ), .QN(n9336));
   SDFFARX1 \key_mem_reg[4][65]  (.D(n4360), .SI(n9209), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[4][65] ), .QN(n9208));
   SDFFARX1 \key_mem_reg[5][65]  (.D(n4361), .SI(n9082), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[5][65] ), .QN(n9081));
   SDFFARX1 \key_mem_reg[6][65]  (.D(n4362), .SI(n8954), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[6][65] ), .QN(n8953));
   SDFFARX1 \key_mem_reg[7][65]  (.D(n4363), .SI(n8826), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[7][65] ), .QN(n8825));
   SDFFARX1 \key_mem_reg[8][65]  (.D(n4364), .SI(n8698), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[8][65] ), .QN(n8697));
   SDFFARX1 \key_mem_reg[9][65]  (.D(n4365), .SI(n8570), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[9][65] ), .QN(n8569));
   SDFFARX1 \key_mem_reg[10][65]  (.D(n4366), .SI(n8442), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[10][65] ), .QN(n8441));
   SDFFARX1 \key_mem_reg[11][65]  (.D(n4367), .SI(n8314), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[11][65] ), .QN(n8313));
   SDFFARX1 \key_mem_reg[12][65]  (.D(n4368), .SI(n8187), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[12][65] ), .QN(n8186));
   SDFFARX1 \key_mem_reg[13][65]  (.D(n4369), .SI(n8059), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[13][65] ), .QN(n8058));
   SDFFARX1 \key_mem_reg[14][65]  (.D(n4370), .SI(n7931), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(\key_mem[14][65] ), .QN(n7930));
   SDFFARX1 \prev_key1_reg_reg[64]  (.D(n5409), .SI(n7693), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7405), .Q(prev_key1_reg[64]), .QN(n7692));
   SDFFARX1 \prev_key0_reg_reg[64]  (.D(n5536), .SI(n7804), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(prev_key0_reg[64]), .QN(n7803));
   SDFFARX1 \key_mem_reg[0][64]  (.D(n4371), .SI(n9722), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[0][64] ), .QN(n9721));
   SDFFARX1 \key_mem_reg[1][64]  (.D(n4372), .SI(n9594), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[1][64] ), .QN(n9593));
   SDFFARX1 \key_mem_reg[2][64]  (.D(n4373), .SI(n9466), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[2][64] ), .QN(n9465));
   SDFFARX1 \key_mem_reg[3][64]  (.D(n4374), .SI(n9338), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[3][64] ), .QN(n9337));
   SDFFARX1 \key_mem_reg[4][64]  (.D(n4375), .SI(n9210), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[4][64] ), .QN(n9209));
   SDFFARX1 \key_mem_reg[5][64]  (.D(n4376), .SI(n9083), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[5][64] ), .QN(n9082));
   SDFFARX1 \key_mem_reg[6][64]  (.D(n4377), .SI(n8955), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[6][64] ), .QN(n8954));
   SDFFARX1 \key_mem_reg[7][64]  (.D(n4378), .SI(n8827), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[7][64] ), .QN(n8826));
   SDFFARX1 \key_mem_reg[8][64]  (.D(n4379), .SI(n8699), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[8][64] ), .QN(n8698));
   SDFFARX1 \key_mem_reg[9][64]  (.D(n4380), .SI(n8571), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[9][64] ), .QN(n8570));
   SDFFARX1 \key_mem_reg[10][64]  (.D(n4381), .SI(n8443), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7404), .Q(\key_mem[10][64] ), .QN(n8442));
   SDFFARX1 \key_mem_reg[11][64]  (.D(n4382), .SI(n8315), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[11][64] ), .QN(n8314));
   SDFFARX1 \key_mem_reg[12][64]  (.D(n4383), .SI(n8188), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[12][64] ), .QN(n8187));
   SDFFARX1 \key_mem_reg[13][64]  (.D(n4384), .SI(n8060), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[13][64] ), .QN(n8059));
   SDFFARX1 \key_mem_reg[14][64]  (.D(n4385), .SI(n7932), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[14][64] ), .QN(n7931));
   SDFFARX1 \prev_key1_reg_reg[63]  (.D(n5410), .SI(n7694), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(prev_key1_reg[63]), .QN(n7693));
   SDFFARX1 \prev_key0_reg_reg[63]  (.D(n5537), .SI(n7805), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(prev_key0_reg[63]), .QN(n7804));
   SDFFARX1 \key_mem_reg[0][63]  (.D(n4386), .SI(n9723), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[0][63] ), .QN(n9722));
   SDFFARX1 \key_mem_reg[1][63]  (.D(n4387), .SI(n9595), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[1][63] ), .QN(n9594));
   SDFFARX1 \key_mem_reg[2][63]  (.D(n4388), .SI(n9467), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[2][63] ), .QN(n9466));
   SDFFARX1 \key_mem_reg[3][63]  (.D(n4389), .SI(n9339), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[3][63] ), .QN(n9338));
   SDFFARX1 \key_mem_reg[4][63]  (.D(n4390), .SI(n9211), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[4][63] ), .QN(n9210));
   SDFFARX1 \key_mem_reg[5][63]  (.D(n4391), .SI(n9084), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7403), .Q(\key_mem[5][63] ), .QN(n9083));
   SDFFARX1 \key_mem_reg[6][63]  (.D(n4392), .SI(n8956), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[6][63] ), .QN(n8955));
   SDFFARX1 \key_mem_reg[7][63]  (.D(n4393), .SI(n8828), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[7][63] ), .QN(n8827));
   SDFFARX1 \key_mem_reg[8][63]  (.D(n4394), .SI(n8700), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[8][63] ), .QN(n8699));
   SDFFARX1 \key_mem_reg[9][63]  (.D(n4395), .SI(n8572), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[9][63] ), .QN(n8571));
   SDFFARX1 \key_mem_reg[10][63]  (.D(n4396), .SI(n8444), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[10][63] ), .QN(n8443));
   SDFFARX1 \key_mem_reg[11][63]  (.D(n4397), .SI(n8316), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[11][63] ), .QN(n8315));
   SDFFARX1 \key_mem_reg[12][63]  (.D(n4398), .SI(n8189), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[12][63] ), .QN(n8188));
   SDFFARX1 \key_mem_reg[13][63]  (.D(n4399), .SI(n8061), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[13][63] ), .QN(n8060));
   SDFFARX1 \key_mem_reg[14][63]  (.D(n4400), .SI(n7933), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[14][63] ), .QN(n7932));
   SDFFARX1 \prev_key1_reg_reg[62]  (.D(n5411), .SI(n7695), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(prev_key1_reg[62]), .QN(n7694));
   SDFFARX1 \prev_key0_reg_reg[62]  (.D(n5538), .SI(n7806), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(prev_key0_reg[62]), .QN(n7805));
   SDFFARX1 \key_mem_reg[0][62]  (.D(n4401), .SI(n9724), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7402), .Q(\key_mem[0][62] ), .QN(n9723));
   SDFFARX1 \key_mem_reg[1][62]  (.D(n4402), .SI(n9596), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[1][62] ), .QN(n9595));
   SDFFARX1 \key_mem_reg[2][62]  (.D(n4403), .SI(n9468), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[2][62] ), .QN(n9467));
   SDFFARX1 \key_mem_reg[3][62]  (.D(n4404), .SI(n9340), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[3][62] ), .QN(n9339));
   SDFFARX1 \key_mem_reg[4][62]  (.D(n4405), .SI(n9212), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[4][62] ), .QN(n9211));
   SDFFARX1 \key_mem_reg[5][62]  (.D(n4406), .SI(n9085), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[5][62] ), .QN(n9084));
   SDFFARX1 \key_mem_reg[6][62]  (.D(n4407), .SI(n8957), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[6][62] ), .QN(n8956));
   SDFFARX1 \key_mem_reg[7][62]  (.D(n4408), .SI(n8829), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[7][62] ), .QN(n8828));
   SDFFARX1 \key_mem_reg[8][62]  (.D(n4409), .SI(n8701), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[8][62] ), .QN(n8700));
   SDFFARX1 \key_mem_reg[9][62]  (.D(n4410), .SI(n8573), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[9][62] ), .QN(n8572));
   SDFFARX1 \key_mem_reg[10][62]  (.D(n4411), .SI(n8445), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[10][62] ), .QN(n8444));
   SDFFARX1 \key_mem_reg[11][62]  (.D(n4412), .SI(n8317), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[11][62] ), .QN(n8316));
   SDFFARX1 \key_mem_reg[12][62]  (.D(n4413), .SI(n8190), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7401), .Q(\key_mem[12][62] ), .QN(n8189));
   SDFFARX1 \key_mem_reg[13][62]  (.D(n4414), .SI(n8062), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[13][62] ), .QN(n8061));
   SDFFARX1 \key_mem_reg[14][62]  (.D(n4415), .SI(n7934), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[14][62] ), .QN(n7933));
   SDFFARX1 \prev_key1_reg_reg[61]  (.D(n5412), .SI(n7696), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(prev_key1_reg[61]), .QN(n7695));
   SDFFARX1 \prev_key0_reg_reg[61]  (.D(n5539), .SI(n7807), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(prev_key0_reg[61]), .QN(n7806));
   SDFFARX1 \key_mem_reg[0][61]  (.D(n4416), .SI(n9725), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[0][61] ), .QN(n9724));
   SDFFARX1 \key_mem_reg[1][61]  (.D(n4417), .SI(n9597), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[1][61] ), .QN(n9596));
   SDFFARX1 \key_mem_reg[2][61]  (.D(n4418), .SI(n9469), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[2][61] ), .QN(n9468));
   SDFFARX1 \key_mem_reg[3][61]  (.D(n4419), .SI(n9341), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[3][61] ), .QN(n9340));
   SDFFARX1 \key_mem_reg[4][61]  (.D(n4420), .SI(n9213), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[4][61] ), .QN(n9212));
   SDFFARX1 \key_mem_reg[5][61]  (.D(n4421), .SI(n9086), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[5][61] ), .QN(n9085));
   SDFFARX1 \key_mem_reg[6][61]  (.D(n4422), .SI(n8958), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[6][61] ), .QN(n8957));
   SDFFARX1 \key_mem_reg[7][61]  (.D(n4423), .SI(n8830), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7400), .Q(\key_mem[7][61] ), .QN(n8829));
   SDFFARX1 \key_mem_reg[8][61]  (.D(n4424), .SI(n8702), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[8][61] ), .QN(n8701));
   SDFFARX1 \key_mem_reg[9][61]  (.D(n4425), .SI(n8574), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[9][61] ), .QN(n8573));
   SDFFARX1 \key_mem_reg[10][61]  (.D(n4426), .SI(n8446), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[10][61] ), .QN(n8445));
   SDFFARX1 \key_mem_reg[11][61]  (.D(n4427), .SI(n8318), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[11][61] ), .QN(n8317));
   SDFFARX1 \key_mem_reg[12][61]  (.D(n4428), .SI(n8191), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[12][61] ), .QN(n8190));
   SDFFARX1 \key_mem_reg[13][61]  (.D(n4429), .SI(n8063), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[13][61] ), .QN(n8062));
   SDFFARX1 \key_mem_reg[14][61]  (.D(n4430), .SI(n7935), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[14][61] ), .QN(n7934));
   SDFFARX1 \prev_key1_reg_reg[60]  (.D(n5413), .SI(n7697), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(prev_key1_reg[60]), .QN(n7696));
   SDFFARX1 \prev_key0_reg_reg[60]  (.D(n5540), .SI(n7808), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(prev_key0_reg[60]), .QN(n7807));
   SDFFARX1 \key_mem_reg[0][60]  (.D(n4431), .SI(n9726), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[0][60] ), .QN(n9725));
   SDFFARX1 \key_mem_reg[1][60]  (.D(n4432), .SI(n9598), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[1][60] ), .QN(n9597));
   SDFFARX1 \key_mem_reg[2][60]  (.D(n4433), .SI(n9470), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7399), .Q(\key_mem[2][60] ), .QN(n9469));
   SDFFARX1 \key_mem_reg[3][60]  (.D(n4434), .SI(n9342), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[3][60] ), .QN(n9341));
   SDFFARX1 \key_mem_reg[4][60]  (.D(n4435), .SI(n9214), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[4][60] ), .QN(n9213));
   SDFFARX1 \key_mem_reg[5][60]  (.D(n4436), .SI(n9087), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[5][60] ), .QN(n9086));
   SDFFARX1 \key_mem_reg[6][60]  (.D(n4437), .SI(n8959), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[6][60] ), .QN(n8958));
   SDFFARX1 \key_mem_reg[7][60]  (.D(n4438), .SI(n8831), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[7][60] ), .QN(n8830));
   SDFFARX1 \key_mem_reg[8][60]  (.D(n4439), .SI(n8703), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[8][60] ), .QN(n8702));
   SDFFARX1 \key_mem_reg[9][60]  (.D(n4440), .SI(n8575), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[9][60] ), .QN(n8574));
   SDFFARX1 \key_mem_reg[10][60]  (.D(n4441), .SI(n8447), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[10][60] ), .QN(n8446));
   SDFFARX1 \key_mem_reg[11][60]  (.D(n4442), .SI(n8319), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[11][60] ), .QN(n8318));
   SDFFARX1 \key_mem_reg[12][60]  (.D(n4443), .SI(n8192), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[12][60] ), .QN(n8191));
   SDFFARX1 \key_mem_reg[13][60]  (.D(n4444), .SI(n8064), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[13][60] ), .QN(n8063));
   SDFFARX1 \key_mem_reg[14][60]  (.D(n4445), .SI(n7936), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7398), .Q(\key_mem[14][60] ), .QN(n7935));
   SDFFARX1 \prev_key1_reg_reg[59]  (.D(n5414), .SI(n7698), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(prev_key1_reg[59]), .QN(n7697));
   SDFFARX1 \prev_key0_reg_reg[59]  (.D(n5541), .SI(n7809), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(prev_key0_reg[59]), .QN(n7808));
   SDFFARX1 \key_mem_reg[0][59]  (.D(n4446), .SI(n9727), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[0][59] ), .QN(n9726));
   SDFFARX1 \key_mem_reg[1][59]  (.D(n4447), .SI(n9599), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[1][59] ), .QN(n9598));
   SDFFARX1 \key_mem_reg[2][59]  (.D(n4448), .SI(n9471), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[2][59] ), .QN(n9470));
   SDFFARX1 \key_mem_reg[3][59]  (.D(n4449), .SI(n9343), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[3][59] ), .QN(n9342));
   SDFFARX1 \key_mem_reg[4][59]  (.D(n4450), .SI(n9215), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[4][59] ), .QN(n9214));
   SDFFARX1 \key_mem_reg[5][59]  (.D(n4451), .SI(n9088), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[5][59] ), .QN(n9087));
   SDFFARX1 \key_mem_reg[6][59]  (.D(n4452), .SI(n8960), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[6][59] ), .QN(n8959));
   SDFFARX1 \key_mem_reg[7][59]  (.D(n4453), .SI(n8832), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[7][59] ), .QN(n8831));
   SDFFARX1 \key_mem_reg[8][59]  (.D(n4454), .SI(n8704), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[8][59] ), .QN(n8703));
   SDFFARX1 \key_mem_reg[9][59]  (.D(n4455), .SI(n8576), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7397), .Q(\key_mem[9][59] ), .QN(n8575));
   SDFFARX1 \key_mem_reg[10][59]  (.D(n4456), .SI(n8448), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[10][59] ), .QN(n8447));
   SDFFARX1 \key_mem_reg[11][59]  (.D(n4457), .SI(n8320), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[11][59] ), .QN(n8319));
   SDFFARX1 \key_mem_reg[12][59]  (.D(n4458), .SI(n8193), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[12][59] ), .QN(n8192));
   SDFFARX1 \key_mem_reg[13][59]  (.D(n4459), .SI(n8065), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[13][59] ), .QN(n8064));
   SDFFARX1 \key_mem_reg[14][59]  (.D(n4460), .SI(n7937), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[14][59] ), .QN(n7936));
   SDFFARX1 \prev_key1_reg_reg[58]  (.D(n5415), .SI(n7699), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(prev_key1_reg[58]), .QN(n7698));
   SDFFARX1 \prev_key0_reg_reg[58]  (.D(n5542), .SI(n7810), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(prev_key0_reg[58]), .QN(n7809));
   SDFFARX1 \key_mem_reg[0][58]  (.D(n4461), .SI(n9728), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[0][58] ), .QN(n9727));
   SDFFARX1 \key_mem_reg[1][58]  (.D(n4462), .SI(n9600), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[1][58] ), .QN(n9599));
   SDFFARX1 \key_mem_reg[2][58]  (.D(n4463), .SI(n9472), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[2][58] ), .QN(n9471));
   SDFFARX1 \key_mem_reg[3][58]  (.D(n4464), .SI(n9344), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[3][58] ), .QN(n9343));
   SDFFARX1 \key_mem_reg[4][58]  (.D(n4465), .SI(n9216), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7396), .Q(\key_mem[4][58] ), .QN(n9215));
   SDFFARX1 \key_mem_reg[5][58]  (.D(n4466), .SI(n9089), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[5][58] ), .QN(n9088));
   SDFFARX1 \key_mem_reg[6][58]  (.D(n4467), .SI(n8961), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[6][58] ), .QN(n8960));
   SDFFARX1 \key_mem_reg[7][58]  (.D(n4468), .SI(n8833), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[7][58] ), .QN(n8832));
   SDFFARX1 \key_mem_reg[8][58]  (.D(n4469), .SI(n8705), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[8][58] ), .QN(n8704));
   SDFFARX1 \key_mem_reg[9][58]  (.D(n4470), .SI(n8577), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[9][58] ), .QN(n8576));
   SDFFARX1 \key_mem_reg[10][58]  (.D(n4471), .SI(n8449), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[10][58] ), .QN(n8448));
   SDFFARX1 \key_mem_reg[11][58]  (.D(n4472), .SI(n8321), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[11][58] ), .QN(n8320));
   SDFFARX1 \key_mem_reg[12][58]  (.D(n4473), .SI(n8194), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[12][58] ), .QN(n8193));
   SDFFARX1 \key_mem_reg[13][58]  (.D(n4474), .SI(n8066), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[13][58] ), .QN(n8065));
   SDFFARX1 \key_mem_reg[14][58]  (.D(n4475), .SI(n7938), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(\key_mem[14][58] ), .QN(n7937));
   SDFFARX1 \prev_key1_reg_reg[57]  (.D(n5416), .SI(n1), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(prev_key1_reg[57]), .QN(n7699));
   SDFFARX1 \prev_key0_reg_reg[57]  (.D(n5543), .SI(n7811), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7395), .Q(prev_key0_reg[57]), .QN(n7810));
   SDFFARX1 \key_mem_reg[0][57]  (.D(n4476), .SI(n9729), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[0][57] ), .QN(n9728));
   SDFFARX1 \key_mem_reg[1][57]  (.D(n4477), .SI(n9601), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[1][57] ), .QN(n9600));
   SDFFARX1 \key_mem_reg[2][57]  (.D(n4478), .SI(n9473), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[2][57] ), .QN(n9472));
   SDFFARX1 \key_mem_reg[3][57]  (.D(n4479), .SI(n9345), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[3][57] ), .QN(n9344));
   SDFFARX1 \key_mem_reg[4][57]  (.D(n4480), .SI(n9217), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[4][57] ), .QN(n9216));
   SDFFARX1 \key_mem_reg[5][57]  (.D(n4481), .SI(n9090), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[5][57] ), .QN(n9089));
   SDFFARX1 \key_mem_reg[6][57]  (.D(n4482), .SI(n8962), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[6][57] ), .QN(n8961));
   SDFFARX1 \key_mem_reg[7][57]  (.D(n4483), .SI(n8834), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[7][57] ), .QN(n8833));
   SDFFARX1 \key_mem_reg[8][57]  (.D(n4484), .SI(n8706), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[8][57] ), .QN(n8705));
   SDFFARX1 \key_mem_reg[9][57]  (.D(n4485), .SI(n8578), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[9][57] ), .QN(n8577));
   SDFFARX1 \key_mem_reg[10][57]  (.D(n4486), .SI(n8450), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[10][57] ), .QN(n8449));
   SDFFARX1 \key_mem_reg[11][57]  (.D(n4487), .SI(n8322), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7394), .Q(\key_mem[11][57] ), .QN(n8321));
   SDFFARX1 \key_mem_reg[12][57]  (.D(n4488), .SI(n8195), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[12][57] ), .QN(n8194));
   SDFFARX1 \key_mem_reg[13][57]  (.D(n4489), .SI(n8067), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[13][57] ), .QN(n8066));
   SDFFARX1 \key_mem_reg[14][57]  (.D(n4490), .SI(n7939), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[14][57] ), .QN(n7938));
   SDFFARX1 \prev_key1_reg_reg[56]  (.D(n5417), .SI(n7700), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(prev_key1_reg[56]), .QN(n1));
   SDFFARX1 \prev_key0_reg_reg[56]  (.D(n5544), .SI(n7812), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(prev_key0_reg[56]), .QN(n7811));
   SDFFARX1 \key_mem_reg[0][56]  (.D(n4491), .SI(n9730), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[0][56] ), .QN(n9729));
   SDFFARX1 \key_mem_reg[1][56]  (.D(n4492), .SI(n9602), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[1][56] ), .QN(n9601));
   SDFFARX1 \key_mem_reg[2][56]  (.D(n4493), .SI(n9474), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[2][56] ), .QN(n9473));
   SDFFARX1 \key_mem_reg[3][56]  (.D(n4494), .SI(n9346), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[3][56] ), .QN(n9345));
   SDFFARX1 \key_mem_reg[4][56]  (.D(n4495), .SI(n9218), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[4][56] ), .QN(n9217));
   SDFFARX1 \key_mem_reg[5][56]  (.D(n4496), .SI(n9091), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[5][56] ), .QN(n9090));
   SDFFARX1 \key_mem_reg[6][56]  (.D(n4497), .SI(n8963), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7393), .Q(\key_mem[6][56] ), .QN(n8962));
   SDFFARX1 \key_mem_reg[7][56]  (.D(n4498), .SI(n8835), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[7][56] ), .QN(n8834));
   SDFFARX1 \key_mem_reg[8][56]  (.D(n4499), .SI(n8707), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[8][56] ), .QN(n8706));
   SDFFARX1 \key_mem_reg[9][56]  (.D(n4500), .SI(n8579), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[9][56] ), .QN(n8578));
   SDFFARX1 \key_mem_reg[10][56]  (.D(n4501), .SI(n8451), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[10][56] ), .QN(n8450));
   SDFFARX1 \key_mem_reg[11][56]  (.D(n4502), .SI(n8323), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[11][56] ), .QN(n8322));
   SDFFARX1 \key_mem_reg[12][56]  (.D(n4503), .SI(n8196), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[12][56] ), .QN(n8195));
   SDFFARX1 \key_mem_reg[13][56]  (.D(n4504), .SI(n8068), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[13][56] ), .QN(n8067));
   SDFFARX1 \key_mem_reg[14][56]  (.D(n4505), .SI(n7940), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[14][56] ), .QN(n7939));
   SDFFARX1 \prev_key1_reg_reg[55]  (.D(n5418), .SI(n7701), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(prev_key1_reg[55]), .QN(n7700));
   SDFFARX1 \prev_key0_reg_reg[55]  (.D(n5545), .SI(n7813), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(prev_key0_reg[55]), .QN(n7812));
   SDFFARX1 \key_mem_reg[0][55]  (.D(n4506), .SI(n9731), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[0][55] ), .QN(n9730));
   SDFFARX1 \key_mem_reg[1][55]  (.D(n4507), .SI(n9603), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7392), .Q(\key_mem[1][55] ), .QN(n9602));
   SDFFARX1 \key_mem_reg[2][55]  (.D(n4508), .SI(n9475), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[2][55] ), .QN(n9474));
   SDFFARX1 \key_mem_reg[3][55]  (.D(n4509), .SI(n9347), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[3][55] ), .QN(n9346));
   SDFFARX1 \key_mem_reg[4][55]  (.D(n4510), .SI(n9219), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[4][55] ), .QN(n9218));
   SDFFARX1 \key_mem_reg[5][55]  (.D(n4511), .SI(n9092), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[5][55] ), .QN(n9091));
   SDFFARX1 \key_mem_reg[6][55]  (.D(n4512), .SI(n8964), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[6][55] ), .QN(n8963));
   SDFFARX1 \key_mem_reg[7][55]  (.D(n4513), .SI(n8836), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[7][55] ), .QN(n8835));
   SDFFARX1 \key_mem_reg[8][55]  (.D(n4514), .SI(n8708), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[8][55] ), .QN(n8707));
   SDFFARX1 \key_mem_reg[9][55]  (.D(n4515), .SI(n8580), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[9][55] ), .QN(n8579));
   SDFFARX1 \key_mem_reg[10][55]  (.D(n4516), .SI(n8452), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[10][55] ), .QN(n8451));
   SDFFARX1 \key_mem_reg[11][55]  (.D(n4517), .SI(n8324), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[11][55] ), .QN(n8323));
   SDFFARX1 \key_mem_reg[12][55]  (.D(n4518), .SI(n8197), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[12][55] ), .QN(n8196));
   SDFFARX1 \key_mem_reg[13][55]  (.D(n4519), .SI(n8069), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7391), .Q(\key_mem[13][55] ), .QN(n8068));
   SDFFARX1 \key_mem_reg[14][55]  (.D(n4520), .SI(n7941), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[14][55] ), .QN(n7940));
   SDFFARX1 \prev_key1_reg_reg[54]  (.D(n5419), .SI(n7702), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(prev_key1_reg[54]), .QN(n7701));
   SDFFARX1 \prev_key0_reg_reg[54]  (.D(n5546), .SI(n7814), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(prev_key0_reg[54]), .QN(n7813));
   SDFFARX1 \key_mem_reg[0][54]  (.D(n4521), .SI(n9732), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[0][54] ), .QN(n9731));
   SDFFARX1 \key_mem_reg[1][54]  (.D(n4522), .SI(n9604), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[1][54] ), .QN(n9603));
   SDFFARX1 \key_mem_reg[2][54]  (.D(n4523), .SI(n9476), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[2][54] ), .QN(n9475));
   SDFFARX1 \key_mem_reg[3][54]  (.D(n4524), .SI(n9348), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[3][54] ), .QN(n9347));
   SDFFARX1 \key_mem_reg[4][54]  (.D(n4525), .SI(n9220), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[4][54] ), .QN(n9219));
   SDFFARX1 \key_mem_reg[5][54]  (.D(n4526), .SI(n9093), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[5][54] ), .QN(n9092));
   SDFFARX1 \key_mem_reg[6][54]  (.D(n4527), .SI(n8965), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[6][54] ), .QN(n8964));
   SDFFARX1 \key_mem_reg[7][54]  (.D(n4528), .SI(n8837), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[7][54] ), .QN(n8836));
   SDFFARX1 \key_mem_reg[8][54]  (.D(n4529), .SI(n8709), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7390), .Q(\key_mem[8][54] ), .QN(n8708));
   SDFFARX1 \key_mem_reg[9][54]  (.D(n4530), .SI(n8581), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[9][54] ), .QN(n8580));
   SDFFARX1 \key_mem_reg[10][54]  (.D(n4531), .SI(n8453), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[10][54] ), .QN(n8452));
   SDFFARX1 \key_mem_reg[11][54]  (.D(n4532), .SI(n8325), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[11][54] ), .QN(n8324));
   SDFFARX1 \key_mem_reg[12][54]  (.D(n4533), .SI(n8198), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[12][54] ), .QN(n8197));
   SDFFARX1 \key_mem_reg[13][54]  (.D(n4534), .SI(n8070), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[13][54] ), .QN(n8069));
   SDFFARX1 \key_mem_reg[14][54]  (.D(n4535), .SI(n7942), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[14][54] ), .QN(n7941));
   SDFFARX1 \prev_key1_reg_reg[53]  (.D(n5420), .SI(n7703), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(prev_key1_reg[53]), .QN(n7702));
   SDFFARX1 \prev_key0_reg_reg[53]  (.D(n5547), .SI(n7815), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(prev_key0_reg[53]), .QN(n7814));
   SDFFARX1 \key_mem_reg[0][53]  (.D(n4536), .SI(n9733), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[0][53] ), .QN(n9732));
   SDFFARX1 \key_mem_reg[1][53]  (.D(n4537), .SI(n9605), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[1][53] ), .QN(n9604));
   SDFFARX1 \key_mem_reg[2][53]  (.D(n4538), .SI(n9477), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[2][53] ), .QN(n9476));
   SDFFARX1 \key_mem_reg[3][53]  (.D(n4539), .SI(n9349), .SE(test_se_buf_net3), .CLK(
          clk_buf_net3), .RSTB(n7389), .Q(\key_mem[3][53] ), .QN(n9348));
   SDFFARX1 \key_mem_reg[4][53]  (.D(n4540), .SI(n9221), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[4][53] ), .QN(n9220));
   SDFFARX1 \key_mem_reg[5][53]  (.D(n4541), .SI(n9094), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[5][53] ), .QN(n9093));
   SDFFARX1 \key_mem_reg[6][53]  (.D(n4542), .SI(n8966), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[6][53] ), .QN(n8965));
   SDFFARX1 \key_mem_reg[7][53]  (.D(n4543), .SI(n8838), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[7][53] ), .QN(n8837));
   SDFFARX1 \key_mem_reg[8][53]  (.D(n4544), .SI(n8710), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[8][53] ), .QN(n8709));
   SDFFARX1 \key_mem_reg[9][53]  (.D(n4545), .SI(n8582), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[9][53] ), .QN(n8581));
   SDFFARX1 \key_mem_reg[10][53]  (.D(n4546), .SI(n8454), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[10][53] ), .QN(n8453));
   SDFFARX1 \key_mem_reg[11][53]  (.D(n4547), .SI(n8326), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[11][53] ), .QN(n8325));
   SDFFARX1 \key_mem_reg[12][53]  (.D(n4548), .SI(n8199), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[12][53] ), .QN(n8198));
   SDFFARX1 \key_mem_reg[13][53]  (.D(n4549), .SI(n8071), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[13][53] ), .QN(n8070));
   SDFFARX1 \key_mem_reg[14][53]  (.D(n4550), .SI(n7943), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(\key_mem[14][53] ), .QN(n7942));
   SDFFARX1 \prev_key1_reg_reg[52]  (.D(n5421), .SI(n7704), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7388), .Q(prev_key1_reg[52]), .QN(n7703));
   SDFFARX1 \prev_key0_reg_reg[52]  (.D(n5548), .SI(n7816), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(prev_key0_reg[52]), .QN(n7815));
   SDFFARX1 \key_mem_reg[0][52]  (.D(n4551), .SI(n9734), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[0][52] ), .QN(n9733));
   SDFFARX1 \key_mem_reg[1][52]  (.D(n4552), .SI(n9606), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[1][52] ), .QN(n9605));
   SDFFARX1 \key_mem_reg[2][52]  (.D(n4553), .SI(n9478), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[2][52] ), .QN(n9477));
   SDFFARX1 \key_mem_reg[3][52]  (.D(n4554), .SI(n9350), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[3][52] ), .QN(n9349));
   SDFFARX1 \key_mem_reg[4][52]  (.D(n4555), .SI(n9222), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[4][52] ), .QN(n9221));
   SDFFARX1 \key_mem_reg[5][52]  (.D(n4556), .SI(n9095), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[5][52] ), .QN(n9094));
   SDFFARX1 \key_mem_reg[6][52]  (.D(n4557), .SI(n8967), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[6][52] ), .QN(n8966));
   SDFFARX1 \key_mem_reg[7][52]  (.D(n4558), .SI(n8839), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[7][52] ), .QN(n8838));
   SDFFARX1 \key_mem_reg[8][52]  (.D(n4559), .SI(n8711), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[8][52] ), .QN(n8710));
   SDFFARX1 \key_mem_reg[9][52]  (.D(n4560), .SI(n8583), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[9][52] ), .QN(n8582));
   SDFFARX1 \key_mem_reg[10][52]  (.D(n4561), .SI(n8455), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7387), .Q(\key_mem[10][52] ), .QN(n8454));
   SDFFARX1 \key_mem_reg[11][52]  (.D(n4562), .SI(n8327), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[11][52] ), .QN(n8326));
   SDFFARX1 \key_mem_reg[12][52]  (.D(n4563), .SI(n8200), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[12][52] ), .QN(n8199));
   SDFFARX1 \key_mem_reg[13][52]  (.D(n4564), .SI(n8072), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[13][52] ), .QN(n8071));
   SDFFARX1 \key_mem_reg[14][52]  (.D(n4565), .SI(n7944), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[14][52] ), .QN(n7943));
   SDFFARX1 \prev_key1_reg_reg[51]  (.D(n5422), .SI(n7705), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(prev_key1_reg[51]), .QN(n7704));
   SDFFARX1 \prev_key0_reg_reg[51]  (.D(n5549), .SI(n7817), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(prev_key0_reg[51]), .QN(n7816));
   SDFFARX1 \key_mem_reg[0][51]  (.D(n4566), .SI(n9735), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[0][51] ), .QN(n9734));
   SDFFARX1 \key_mem_reg[1][51]  (.D(n4567), .SI(n9607), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[1][51] ), .QN(n9606));
   SDFFARX1 \key_mem_reg[2][51]  (.D(n4568), .SI(n9479), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[2][51] ), .QN(n9478));
   SDFFARX1 \key_mem_reg[3][51]  (.D(n4569), .SI(n9351), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[3][51] ), .QN(n9350));
   SDFFARX1 \key_mem_reg[4][51]  (.D(n4570), .SI(n9223), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[4][51] ), .QN(n9222));
   SDFFARX1 \key_mem_reg[5][51]  (.D(n4571), .SI(n9096), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7386), .Q(\key_mem[5][51] ), .QN(n9095));
   SDFFARX1 \key_mem_reg[6][51]  (.D(n4572), .SI(n8968), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[6][51] ), .QN(n8967));
   SDFFARX1 \key_mem_reg[7][51]  (.D(n4573), .SI(n8840), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[7][51] ), .QN(n8839));
   SDFFARX1 \key_mem_reg[8][51]  (.D(n4574), .SI(n8712), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[8][51] ), .QN(n8711));
   SDFFARX1 \key_mem_reg[9][51]  (.D(n4575), .SI(n8584), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[9][51] ), .QN(n8583));
   SDFFARX1 \key_mem_reg[10][51]  (.D(n4576), .SI(n8456), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[10][51] ), .QN(n8455));
   SDFFARX1 \key_mem_reg[11][51]  (.D(n4577), .SI(n8328), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[11][51] ), .QN(n8327));
   SDFFARX1 \key_mem_reg[12][51]  (.D(n4578), .SI(n8201), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[12][51] ), .QN(n8200));
   SDFFARX1 \key_mem_reg[13][51]  (.D(n4579), .SI(n8073), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[13][51] ), .QN(n8072));
   SDFFARX1 \key_mem_reg[14][51]  (.D(n4580), .SI(n7945), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[14][51] ), .QN(n7944));
   SDFFARX1 \prev_key1_reg_reg[50]  (.D(n5423), .SI(n7706), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(prev_key1_reg[50]), .QN(n7705));
   SDFFARX1 \prev_key0_reg_reg[50]  (.D(n5550), .SI(n7818), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(prev_key0_reg[50]), .QN(n7817));
   SDFFARX1 \key_mem_reg[0][50]  (.D(n4581), .SI(n9736), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7385), .Q(\key_mem[0][50] ), .QN(n9735));
   SDFFARX1 \key_mem_reg[1][50]  (.D(n4582), .SI(n9608), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[1][50] ), .QN(n9607));
   SDFFARX1 \key_mem_reg[2][50]  (.D(n4583), .SI(n9480), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[2][50] ), .QN(n9479));
   SDFFARX1 \key_mem_reg[3][50]  (.D(n4584), .SI(n9352), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[3][50] ), .QN(n9351));
   SDFFARX1 \key_mem_reg[4][50]  (.D(n4585), .SI(n9224), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[4][50] ), .QN(n9223));
   SDFFARX1 \key_mem_reg[5][50]  (.D(n4586), .SI(n9097), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[5][50] ), .QN(n9096));
   SDFFARX1 \key_mem_reg[6][50]  (.D(n4587), .SI(n8969), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[6][50] ), .QN(n8968));
   SDFFARX1 \key_mem_reg[7][50]  (.D(n4588), .SI(n8841), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[7][50] ), .QN(n8840));
   SDFFARX1 \key_mem_reg[8][50]  (.D(n4589), .SI(n8713), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[8][50] ), .QN(n8712));
   SDFFARX1 \key_mem_reg[9][50]  (.D(n4590), .SI(n8585), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[9][50] ), .QN(n8584));
   SDFFARX1 \key_mem_reg[10][50]  (.D(n4591), .SI(n8457), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[10][50] ), .QN(n8456));
   SDFFARX1 \key_mem_reg[11][50]  (.D(n4592), .SI(n8329), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[11][50] ), .QN(n8328));
   SDFFARX1 \key_mem_reg[12][50]  (.D(n4593), .SI(test_si3), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7384), .Q(\key_mem[12][50] ), .QN(n8201));
   SDFFARX1 \key_mem_reg[13][50]  (.D(n4594), .SI(n8074), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[13][50] ), .QN(n8073));
   SDFFARX1 \key_mem_reg[14][50]  (.D(n4595), .SI(n7946), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[14][50] ), .QN(n7945));
   SDFFARX1 \prev_key1_reg_reg[49]  (.D(n5424), .SI(n7707), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(prev_key1_reg[49]), .QN(n7706));
   SDFFARX1 \prev_key0_reg_reg[49]  (.D(n5551), .SI(n7819), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(prev_key0_reg[49]), .QN(n7818));
   SDFFARX1 \key_mem_reg[0][49]  (.D(n4596), .SI(n9737), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[0][49] ), .QN(n9736));
   SDFFARX1 \key_mem_reg[1][49]  (.D(n4597), .SI(n9609), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[1][49] ), .QN(n9608));
   SDFFARX1 \key_mem_reg[2][49]  (.D(n4598), .SI(n9481), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[2][49] ), .QN(n9480));
   SDFFARX1 \key_mem_reg[3][49]  (.D(n4599), .SI(n9353), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[3][49] ), .QN(n9352));
   SDFFARX1 \key_mem_reg[4][49]  (.D(n4600), .SI(n9225), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[4][49] ), .QN(n9224));
   SDFFARX1 \key_mem_reg[5][49]  (.D(n4601), .SI(n9098), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[5][49] ), .QN(n9097));
   SDFFARX1 \key_mem_reg[6][49]  (.D(n4602), .SI(n8970), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[6][49] ), .QN(n8969));
   SDFFARX1 \key_mem_reg[7][49]  (.D(n4603), .SI(n8842), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7383), .Q(\key_mem[7][49] ), .QN(n8841));
   SDFFARX1 \key_mem_reg[8][49]  (.D(n4604), .SI(n8714), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[8][49] ), .QN(n8713));
   SDFFARX1 \key_mem_reg[9][49]  (.D(n4605), .SI(n8586), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[9][49] ), .QN(n8585));
   SDFFARX1 \key_mem_reg[10][49]  (.D(n4606), .SI(n8458), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[10][49] ), .QN(n8457));
   SDFFARX1 \key_mem_reg[11][49]  (.D(n4607), .SI(n8330), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[11][49] ), .QN(n8329));
   SDFFARX1 \key_mem_reg[12][49]  (.D(n4608), .SI(n8202), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[12][49] ));
   SDFFARX1 \key_mem_reg[13][49]  (.D(n4609), .SI(n8075), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[13][49] ), .QN(n8074));
   SDFFARX1 \key_mem_reg[14][49]  (.D(n4610), .SI(n7947), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[14][49] ), .QN(n7946));
   SDFFARX1 \prev_key1_reg_reg[48]  (.D(n5425), .SI(n7708), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(prev_key1_reg[48]), .QN(n7707));
   SDFFARX1 \prev_key0_reg_reg[48]  (.D(n5552), .SI(n7820), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(prev_key0_reg[48]), .QN(n7819));
   SDFFARX1 \key_mem_reg[0][48]  (.D(n4611), .SI(n9738), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[0][48] ), .QN(n9737));
   SDFFARX1 \key_mem_reg[1][48]  (.D(n4612), .SI(n9610), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[1][48] ), .QN(n9609));
   SDFFARX1 \key_mem_reg[2][48]  (.D(n4613), .SI(n9482), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7382), .Q(\key_mem[2][48] ), .QN(n9481));
   SDFFARX1 \key_mem_reg[3][48]  (.D(n4614), .SI(n9354), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[3][48] ), .QN(n9353));
   SDFFARX1 \key_mem_reg[4][48]  (.D(n4615), .SI(n9226), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[4][48] ), .QN(n9225));
   SDFFARX1 \key_mem_reg[5][48]  (.D(n4616), .SI(n9099), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[5][48] ), .QN(n9098));
   SDFFARX1 \key_mem_reg[6][48]  (.D(n4617), .SI(n8971), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[6][48] ), .QN(n8970));
   SDFFARX1 \key_mem_reg[7][48]  (.D(n4618), .SI(n8843), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[7][48] ), .QN(n8842));
   SDFFARX1 \key_mem_reg[8][48]  (.D(n4619), .SI(n8715), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[8][48] ), .QN(n8714));
   SDFFARX1 \key_mem_reg[9][48]  (.D(n4620), .SI(n8587), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[9][48] ), .QN(n8586));
   SDFFARX1 \key_mem_reg[10][48]  (.D(n4621), .SI(n8459), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[10][48] ), .QN(n8458));
   SDFFARX1 \key_mem_reg[11][48]  (.D(n4622), .SI(n8331), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[11][48] ), .QN(n8330));
   SDFFARX1 \key_mem_reg[12][48]  (.D(n4623), .SI(n8203), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[12][48] ), .QN(n8202));
   SDFFARX1 \key_mem_reg[13][48]  (.D(n4624), .SI(n8076), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[13][48] ), .QN(n8075));
   SDFFARX1 \key_mem_reg[14][48]  (.D(n4625), .SI(n7948), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7381), .Q(\key_mem[14][48] ), .QN(n7947));
   SDFFARX1 \prev_key1_reg_reg[47]  (.D(n5426), .SI(n7709), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(prev_key1_reg[47]), .QN(n7708));
   SDFFARX1 \prev_key0_reg_reg[47]  (.D(n5553), .SI(n7821), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(prev_key0_reg[47]), .QN(n7820));
   SDFFARX1 \key_mem_reg[0][47]  (.D(n4626), .SI(n9739), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[0][47] ), .QN(n9738));
   SDFFARX1 \key_mem_reg[1][47]  (.D(n4627), .SI(n9611), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[1][47] ), .QN(n9610));
   SDFFARX1 \key_mem_reg[2][47]  (.D(n4628), .SI(n9483), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[2][47] ), .QN(n9482));
   SDFFARX1 \key_mem_reg[3][47]  (.D(n4629), .SI(n9355), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[3][47] ), .QN(n9354));
   SDFFARX1 \key_mem_reg[4][47]  (.D(n4630), .SI(n9227), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[4][47] ), .QN(n9226));
   SDFFARX1 \key_mem_reg[5][47]  (.D(n4631), .SI(n9100), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[5][47] ), .QN(n9099));
   SDFFARX1 \key_mem_reg[6][47]  (.D(n4632), .SI(n8972), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[6][47] ), .QN(n8971));
   SDFFARX1 \key_mem_reg[7][47]  (.D(n4633), .SI(n8844), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[7][47] ), .QN(n8843));
   SDFFARX1 \key_mem_reg[8][47]  (.D(n4634), .SI(n8716), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[8][47] ), .QN(n8715));
   SDFFARX1 \key_mem_reg[9][47]  (.D(n4635), .SI(n8588), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7380), .Q(\key_mem[9][47] ), .QN(n8587));
   SDFFARX1 \key_mem_reg[10][47]  (.D(n4636), .SI(n8460), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[10][47] ), .QN(n8459));
   SDFFARX1 \key_mem_reg[11][47]  (.D(n4637), .SI(n8332), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[11][47] ), .QN(n8331));
   SDFFARX1 \key_mem_reg[12][47]  (.D(n4638), .SI(n8204), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[12][47] ), .QN(n8203));
   SDFFARX1 \key_mem_reg[13][47]  (.D(n4639), .SI(n8077), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[13][47] ), .QN(n8076));
   SDFFARX1 \key_mem_reg[14][47]  (.D(n4640), .SI(n7949), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[14][47] ), .QN(n7948));
   SDFFARX1 \prev_key1_reg_reg[46]  (.D(n5427), .SI(n7710), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(prev_key1_reg[46]), .QN(n7709));
   SDFFARX1 \prev_key0_reg_reg[46]  (.D(n5554), .SI(n7822), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(prev_key0_reg[46]), .QN(n7821));
   SDFFARX1 \key_mem_reg[0][46]  (.D(n4641), .SI(n9740), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[0][46] ), .QN(n9739));
   SDFFARX1 \key_mem_reg[1][46]  (.D(n4642), .SI(n9612), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[1][46] ), .QN(n9611));
   SDFFARX1 \key_mem_reg[2][46]  (.D(n4643), .SI(n9484), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[2][46] ), .QN(n9483));
   SDFFARX1 \key_mem_reg[3][46]  (.D(n4644), .SI(n9356), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[3][46] ), .QN(n9355));
   SDFFARX1 \key_mem_reg[4][46]  (.D(n4645), .SI(n9228), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7379), .Q(\key_mem[4][46] ), .QN(n9227));
   SDFFARX1 \key_mem_reg[5][46]  (.D(n4646), .SI(n9101), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[5][46] ), .QN(n9100));
   SDFFARX1 \key_mem_reg[6][46]  (.D(n4647), .SI(n8973), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[6][46] ), .QN(n8972));
   SDFFARX1 \key_mem_reg[7][46]  (.D(n4648), .SI(n8845), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[7][46] ), .QN(n8844));
   SDFFARX1 \key_mem_reg[8][46]  (.D(n4649), .SI(n8717), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[8][46] ), .QN(n8716));
   SDFFARX1 \key_mem_reg[9][46]  (.D(n4650), .SI(n8589), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[9][46] ), .QN(n8588));
   SDFFARX1 \key_mem_reg[10][46]  (.D(n4651), .SI(n8461), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[10][46] ), .QN(n8460));
   SDFFARX1 \key_mem_reg[11][46]  (.D(n4652), .SI(n8333), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[11][46] ), .QN(n8332));
   SDFFARX1 \key_mem_reg[12][46]  (.D(n4653), .SI(n8205), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[12][46] ), .QN(n8204));
   SDFFARX1 \key_mem_reg[13][46]  (.D(n4654), .SI(n8078), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[13][46] ), .QN(n8077));
   SDFFARX1 \key_mem_reg[14][46]  (.D(n4655), .SI(n7950), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(\key_mem[14][46] ), .QN(n7949));
   SDFFARX1 \prev_key1_reg_reg[45]  (.D(n5428), .SI(n7711), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(prev_key1_reg[45]), .QN(n7710));
   SDFFARX1 \prev_key0_reg_reg[45]  (.D(n5555), .SI(n7823), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7378), .Q(prev_key0_reg[45]), .QN(n7822));
   SDFFARX1 \key_mem_reg[0][45]  (.D(n4656), .SI(n9741), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[0][45] ), .QN(n9740));
   SDFFARX1 \key_mem_reg[1][45]  (.D(n4657), .SI(n9613), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[1][45] ), .QN(n9612));
   SDFFARX1 \key_mem_reg[2][45]  (.D(n4658), .SI(n9485), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[2][45] ), .QN(n9484));
   SDFFARX1 \key_mem_reg[3][45]  (.D(n4659), .SI(n9357), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[3][45] ), .QN(n9356));
   SDFFARX1 \key_mem_reg[4][45]  (.D(n4660), .SI(n9229), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[4][45] ), .QN(n9228));
   SDFFARX1 \key_mem_reg[5][45]  (.D(n4661), .SI(n9102), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[5][45] ), .QN(n9101));
   SDFFARX1 \key_mem_reg[6][45]  (.D(n4662), .SI(n8974), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[6][45] ), .QN(n8973));
   SDFFARX1 \key_mem_reg[7][45]  (.D(n4663), .SI(n8846), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[7][45] ), .QN(n8845));
   SDFFARX1 \key_mem_reg[8][45]  (.D(n4664), .SI(n8718), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[8][45] ), .QN(n8717));
   SDFFARX1 \key_mem_reg[9][45]  (.D(n4665), .SI(n8590), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[9][45] ), .QN(n8589));
   SDFFARX1 \key_mem_reg[10][45]  (.D(n4666), .SI(n8462), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[10][45] ), .QN(n8461));
   SDFFARX1 \key_mem_reg[11][45]  (.D(n4667), .SI(n8334), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7377), .Q(\key_mem[11][45] ), .QN(n8333));
   SDFFARX1 \key_mem_reg[12][45]  (.D(n4668), .SI(n8206), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[12][45] ), .QN(n8205));
   SDFFARX1 \key_mem_reg[13][45]  (.D(n4669), .SI(n8079), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[13][45] ), .QN(n8078));
   SDFFARX1 \key_mem_reg[14][45]  (.D(n4670), .SI(n7951), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[14][45] ), .QN(n7950));
   SDFFARX1 \prev_key1_reg_reg[44]  (.D(n5429), .SI(n7712), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(prev_key1_reg[44]), .QN(n7711));
   SDFFARX1 \prev_key0_reg_reg[44]  (.D(n5556), .SI(n7824), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(prev_key0_reg[44]), .QN(n7823));
   SDFFARX1 \key_mem_reg[0][44]  (.D(n4671), .SI(n9742), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[0][44] ), .QN(n9741));
   SDFFARX1 \key_mem_reg[1][44]  (.D(n4672), .SI(n9614), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[1][44] ), .QN(n9613));
   SDFFARX1 \key_mem_reg[2][44]  (.D(n4673), .SI(n9486), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[2][44] ), .QN(n9485));
   SDFFARX1 \key_mem_reg[3][44]  (.D(n4674), .SI(n9358), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[3][44] ), .QN(n9357));
   SDFFARX1 \key_mem_reg[4][44]  (.D(n4675), .SI(n9230), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[4][44] ), .QN(n9229));
   SDFFARX1 \key_mem_reg[5][44]  (.D(n4676), .SI(n9103), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[5][44] ), .QN(n9102));
   SDFFARX1 \key_mem_reg[6][44]  (.D(n4677), .SI(n8975), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7376), .Q(\key_mem[6][44] ), .QN(n8974));
   SDFFARX1 \key_mem_reg[7][44]  (.D(n4678), .SI(n8847), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[7][44] ), .QN(n8846));
   SDFFARX1 \key_mem_reg[8][44]  (.D(n4679), .SI(n8719), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[8][44] ), .QN(n8718));
   SDFFARX1 \key_mem_reg[9][44]  (.D(n4680), .SI(n8591), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[9][44] ), .QN(n8590));
   SDFFARX1 \key_mem_reg[10][44]  (.D(n4681), .SI(n8463), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[10][44] ), .QN(n8462));
   SDFFARX1 \key_mem_reg[11][44]  (.D(n4682), .SI(n8335), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[11][44] ), .QN(n8334));
   SDFFARX1 \key_mem_reg[12][44]  (.D(n4683), .SI(n8207), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[12][44] ), .QN(n8206));
   SDFFARX1 \key_mem_reg[13][44]  (.D(n4684), .SI(n8080), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[13][44] ), .QN(n8079));
   SDFFARX1 \key_mem_reg[14][44]  (.D(n4685), .SI(n7952), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[14][44] ), .QN(n7951));
   SDFFARX1 \prev_key1_reg_reg[43]  (.D(n5430), .SI(n7713), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(prev_key1_reg[43]), .QN(n7712));
   SDFFARX1 \prev_key0_reg_reg[43]  (.D(n5557), .SI(n7825), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(prev_key0_reg[43]), .QN(n7824));
   SDFFARX1 \key_mem_reg[0][43]  (.D(n4686), .SI(n9743), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[0][43] ), .QN(n9742));
   SDFFARX1 \key_mem_reg[1][43]  (.D(n4687), .SI(n9615), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7375), .Q(\key_mem[1][43] ), .QN(n9614));
   SDFFARX1 \key_mem_reg[2][43]  (.D(n4688), .SI(n9487), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[2][43] ), .QN(n9486));
   SDFFARX1 \key_mem_reg[3][43]  (.D(n4689), .SI(n9359), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[3][43] ), .QN(n9358));
   SDFFARX1 \key_mem_reg[4][43]  (.D(n4690), .SI(n9231), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[4][43] ), .QN(n9230));
   SDFFARX1 \key_mem_reg[5][43]  (.D(n4691), .SI(n9104), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[5][43] ), .QN(n9103));
   SDFFARX1 \key_mem_reg[6][43]  (.D(n4692), .SI(n8976), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[6][43] ), .QN(n8975));
   SDFFARX1 \key_mem_reg[7][43]  (.D(n4693), .SI(n8848), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[7][43] ), .QN(n8847));
   SDFFARX1 \key_mem_reg[8][43]  (.D(n4694), .SI(n8720), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[8][43] ), .QN(n8719));
   SDFFARX1 \key_mem_reg[9][43]  (.D(n4695), .SI(n8592), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[9][43] ), .QN(n8591));
   SDFFARX1 \key_mem_reg[10][43]  (.D(n4696), .SI(n8464), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[10][43] ), .QN(n8463));
   SDFFARX1 \key_mem_reg[11][43]  (.D(n4697), .SI(n8336), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[11][43] ), .QN(n8335));
   SDFFARX1 \key_mem_reg[12][43]  (.D(n4698), .SI(n8208), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[12][43] ), .QN(n8207));
   SDFFARX1 \key_mem_reg[13][43]  (.D(n4699), .SI(n8081), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7374), .Q(\key_mem[13][43] ), .QN(n8080));
   SDFFARX1 \key_mem_reg[14][43]  (.D(n4700), .SI(n7953), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[14][43] ), .QN(n7952));
   SDFFARX1 \prev_key1_reg_reg[42]  (.D(n5431), .SI(n7714), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(prev_key1_reg[42]), .QN(n7713));
   SDFFARX1 \prev_key0_reg_reg[42]  (.D(n5558), .SI(n7826), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(prev_key0_reg[42]), .QN(n7825));
   SDFFARX1 \key_mem_reg[0][42]  (.D(n4701), .SI(n9744), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[0][42] ), .QN(n9743));
   SDFFARX1 \key_mem_reg[1][42]  (.D(n4702), .SI(n9616), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[1][42] ), .QN(n9615));
   SDFFARX1 \key_mem_reg[2][42]  (.D(n4703), .SI(n9488), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[2][42] ), .QN(n9487));
   SDFFARX1 \key_mem_reg[3][42]  (.D(n4704), .SI(n9360), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[3][42] ), .QN(n9359));
   SDFFARX1 \key_mem_reg[4][42]  (.D(n4705), .SI(n9232), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[4][42] ), .QN(n9231));
   SDFFARX1 \key_mem_reg[5][42]  (.D(n4706), .SI(n9105), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[5][42] ), .QN(n9104));
   SDFFARX1 \key_mem_reg[6][42]  (.D(n4707), .SI(n8977), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[6][42] ), .QN(n8976));
   SDFFARX1 \key_mem_reg[7][42]  (.D(n4708), .SI(n8849), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[7][42] ), .QN(n8848));
   SDFFARX1 \key_mem_reg[8][42]  (.D(n4709), .SI(n8721), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7373), .Q(\key_mem[8][42] ), .QN(n8720));
   SDFFARX1 \key_mem_reg[9][42]  (.D(n4710), .SI(n8593), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[9][42] ), .QN(n8592));
   SDFFARX1 \key_mem_reg[10][42]  (.D(n4711), .SI(n8465), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[10][42] ), .QN(n8464));
   SDFFARX1 \key_mem_reg[11][42]  (.D(n4712), .SI(n8337), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[11][42] ), .QN(n8336));
   SDFFARX1 \key_mem_reg[12][42]  (.D(n4713), .SI(n8209), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[12][42] ), .QN(n8208));
   SDFFARX1 \key_mem_reg[13][42]  (.D(n4714), .SI(n8082), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[13][42] ), .QN(n8081));
   SDFFARX1 \key_mem_reg[14][42]  (.D(n4715), .SI(n7954), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[14][42] ), .QN(n7953));
   SDFFARX1 \prev_key1_reg_reg[41]  (.D(n5432), .SI(n7715), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(prev_key1_reg[41]), .QN(n7714));
   SDFFARX1 \prev_key0_reg_reg[41]  (.D(n5559), .SI(n7827), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(prev_key0_reg[41]), .QN(n7826));
   SDFFARX1 \key_mem_reg[0][41]  (.D(n4716), .SI(n9745), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[0][41] ), .QN(n9744));
   SDFFARX1 \key_mem_reg[1][41]  (.D(n4717), .SI(n9617), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[1][41] ), .QN(n9616));
   SDFFARX1 \key_mem_reg[2][41]  (.D(n4718), .SI(n9489), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[2][41] ), .QN(n9488));
   SDFFARX1 \key_mem_reg[3][41]  (.D(n4719), .SI(n9361), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7372), .Q(\key_mem[3][41] ), .QN(n9360));
   SDFFARX1 \key_mem_reg[4][41]  (.D(n4720), .SI(n9233), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[4][41] ), .QN(n9232));
   SDFFARX1 \key_mem_reg[5][41]  (.D(n4721), .SI(n9106), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[5][41] ), .QN(n9105));
   SDFFARX1 \key_mem_reg[6][41]  (.D(n4722), .SI(n8978), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[6][41] ), .QN(n8977));
   SDFFARX1 \key_mem_reg[7][41]  (.D(n4723), .SI(n8850), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[7][41] ), .QN(n8849));
   SDFFARX1 \key_mem_reg[8][41]  (.D(n4724), .SI(n8722), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[8][41] ), .QN(n8721));
   SDFFARX1 \key_mem_reg[9][41]  (.D(n4725), .SI(n8594), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[9][41] ), .QN(n8593));
   SDFFARX1 \key_mem_reg[10][41]  (.D(n4726), .SI(n8466), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[10][41] ), .QN(n8465));
   SDFFARX1 \key_mem_reg[11][41]  (.D(n4727), .SI(n8338), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[11][41] ), .QN(n8337));
   SDFFARX1 \key_mem_reg[12][41]  (.D(n4728), .SI(n8210), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[12][41] ), .QN(n8209));
   SDFFARX1 \key_mem_reg[13][41]  (.D(n4729), .SI(n8083), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[13][41] ), .QN(n8082));
   SDFFARX1 \key_mem_reg[14][41]  (.D(n4730), .SI(n7955), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(\key_mem[14][41] ), .QN(n7954));
   SDFFARX1 \prev_key1_reg_reg[40]  (.D(n5433), .SI(n7716), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7371), .Q(prev_key1_reg[40]), .QN(n7715));
   SDFFARX1 \prev_key0_reg_reg[40]  (.D(n5560), .SI(n7828), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(prev_key0_reg[40]), .QN(n7827));
   SDFFARX1 \key_mem_reg[0][40]  (.D(n4731), .SI(n9746), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[0][40] ), .QN(n9745));
   SDFFARX1 \key_mem_reg[1][40]  (.D(n4732), .SI(n9618), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[1][40] ), .QN(n9617));
   SDFFARX1 \key_mem_reg[2][40]  (.D(n4733), .SI(n9490), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[2][40] ), .QN(n9489));
   SDFFARX1 \key_mem_reg[3][40]  (.D(n4734), .SI(n9362), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[3][40] ), .QN(n9361));
   SDFFARX1 \key_mem_reg[4][40]  (.D(n4735), .SI(n9234), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[4][40] ), .QN(n9233));
   SDFFARX1 \key_mem_reg[5][40]  (.D(n4736), .SI(n9107), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[5][40] ), .QN(n9106));
   SDFFARX1 \key_mem_reg[6][40]  (.D(n4737), .SI(n8979), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[6][40] ), .QN(n8978));
   SDFFARX1 \key_mem_reg[7][40]  (.D(n4738), .SI(n8851), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[7][40] ), .QN(n8850));
   SDFFARX1 \key_mem_reg[8][40]  (.D(n4739), .SI(n8723), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[8][40] ), .QN(n8722));
   SDFFARX1 \key_mem_reg[9][40]  (.D(n4740), .SI(n8595), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[9][40] ), .QN(n8594));
   SDFFARX1 \key_mem_reg[10][40]  (.D(n4741), .SI(n8467), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7370), .Q(\key_mem[10][40] ), .QN(n8466));
   SDFFARX1 \key_mem_reg[11][40]  (.D(n4742), .SI(n8339), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[11][40] ), .QN(n8338));
   SDFFARX1 \key_mem_reg[12][40]  (.D(n4743), .SI(n8211), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[12][40] ), .QN(n8210));
   SDFFARX1 \key_mem_reg[13][40]  (.D(n4744), .SI(n8084), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[13][40] ), .QN(n8083));
   SDFFARX1 \key_mem_reg[14][40]  (.D(n4745), .SI(n7956), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[14][40] ), .QN(n7955));
   SDFFARX1 \prev_key1_reg_reg[39]  (.D(n5434), .SI(n7717), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(prev_key1_reg[39]), .QN(n7716));
   SDFFARX1 \prev_key0_reg_reg[39]  (.D(n5561), .SI(n7829), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(prev_key0_reg[39]), .QN(n7828));
   SDFFARX1 \key_mem_reg[0][39]  (.D(n4746), .SI(n9747), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[0][39] ), .QN(n9746));
   SDFFARX1 \key_mem_reg[1][39]  (.D(n4747), .SI(n9619), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[1][39] ), .QN(n9618));
   SDFFARX1 \key_mem_reg[2][39]  (.D(n4748), .SI(n9491), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[2][39] ), .QN(n9490));
   SDFFARX1 \key_mem_reg[3][39]  (.D(n4749), .SI(n9363), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[3][39] ), .QN(n9362));
   SDFFARX1 \key_mem_reg[4][39]  (.D(n4750), .SI(n9235), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[4][39] ), .QN(n9234));
   SDFFARX1 \key_mem_reg[5][39]  (.D(n4751), .SI(n9108), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7369), .Q(\key_mem[5][39] ), .QN(n9107));
   SDFFARX1 \key_mem_reg[6][39]  (.D(n4752), .SI(n8980), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[6][39] ), .QN(n8979));
   SDFFARX1 \key_mem_reg[7][39]  (.D(n4753), .SI(n8852), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[7][39] ), .QN(n8851));
   SDFFARX1 \key_mem_reg[8][39]  (.D(n4754), .SI(n8724), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[8][39] ), .QN(n8723));
   SDFFARX1 \key_mem_reg[9][39]  (.D(n4755), .SI(n8596), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[9][39] ), .QN(n8595));
   SDFFARX1 \key_mem_reg[10][39]  (.D(n4756), .SI(n8468), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[10][39] ), .QN(n8467));
   SDFFARX1 \key_mem_reg[11][39]  (.D(n4757), .SI(n8340), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[11][39] ), .QN(n8339));
   SDFFARX1 \key_mem_reg[12][39]  (.D(n4758), .SI(n8212), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[12][39] ), .QN(n8211));
   SDFFARX1 \key_mem_reg[13][39]  (.D(n4759), .SI(n8085), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[13][39] ), .QN(n8084));
   SDFFARX1 \key_mem_reg[14][39]  (.D(n4760), .SI(n7957), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[14][39] ), .QN(n7956));
   SDFFARX1 \prev_key1_reg_reg[38]  (.D(n5435), .SI(n7718), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(prev_key1_reg[38]), .QN(n7717));
   SDFFARX1 \prev_key0_reg_reg[38]  (.D(n5562), .SI(n7830), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(prev_key0_reg[38]), .QN(n7829));
   SDFFARX1 \key_mem_reg[0][38]  (.D(n4761), .SI(n9748), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7368), .Q(\key_mem[0][38] ), .QN(n9747));
   SDFFARX1 \key_mem_reg[1][38]  (.D(n4762), .SI(n9620), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7367), .Q(\key_mem[1][38] ), .QN(n9619));
   SDFFARX1 \key_mem_reg[2][38]  (.D(n4763), .SI(n9492), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7367), .Q(\key_mem[2][38] ), .QN(n9491));
   SDFFARX1 \key_mem_reg[3][38]  (.D(n4764), .SI(n9364), .SE(test_se_buf_net4), .CLK(
          clk_buf_net4), .RSTB(n7367), .Q(\key_mem[3][38] ), .QN(n9363));
   SDFFARX1 \key_mem_reg[4][38]  (.D(n4765), .SI(n9236), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[4][38] ), .QN(n9235));
   SDFFARX1 \key_mem_reg[5][38]  (.D(n4766), .SI(n9109), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[5][38] ), .QN(n9108));
   SDFFARX1 \key_mem_reg[6][38]  (.D(n4767), .SI(n8981), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[6][38] ), .QN(n8980));
   SDFFARX1 \key_mem_reg[7][38]  (.D(n4768), .SI(n8853), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[7][38] ), .QN(n8852));
   SDFFARX1 \key_mem_reg[8][38]  (.D(n4769), .SI(n8725), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[8][38] ), .QN(n8724));
   SDFFARX1 \key_mem_reg[9][38]  (.D(n4770), .SI(n8597), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[9][38] ), .QN(n8596));
   SDFFARX1 \key_mem_reg[10][38]  (.D(n4771), .SI(n8469), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[10][38] ), .QN(n8468));
   SDFFARX1 \key_mem_reg[11][38]  (.D(n4772), .SI(n8341), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[11][38] ), .QN(n8340));
   SDFFARX1 \key_mem_reg[12][38]  (.D(n4773), .SI(n8213), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7367), .Q(\key_mem[12][38] ), .QN(n8212));
   SDFFARX1 \key_mem_reg[13][38]  (.D(n4774), .SI(n8086), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[13][38] ), .QN(n8085));
   SDFFARX1 \key_mem_reg[14][38]  (.D(n4775), .SI(n7958), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[14][38] ), .QN(n7957));
   SDFFARX1 \prev_key1_reg_reg[37]  (.D(n5436), .SI(n7719), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(prev_key1_reg[37]), .QN(n7718));
   SDFFARX1 \prev_key0_reg_reg[37]  (.D(n5563), .SI(n7831), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(prev_key0_reg[37]), .QN(n7830));
   SDFFARX1 \key_mem_reg[0][37]  (.D(n4776), .SI(n9749), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[0][37] ), .QN(n9748));
   SDFFARX1 \key_mem_reg[1][37]  (.D(n4777), .SI(n9621), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[1][37] ), .QN(n9620));
   SDFFARX1 \key_mem_reg[2][37]  (.D(n4778), .SI(n9493), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[2][37] ), .QN(n9492));
   SDFFARX1 \key_mem_reg[3][37]  (.D(n4779), .SI(n9365), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[3][37] ), .QN(n9364));
   SDFFARX1 \key_mem_reg[4][37]  (.D(n4780), .SI(n9237), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[4][37] ), .QN(n9236));
   SDFFARX1 \key_mem_reg[5][37]  (.D(n4781), .SI(n9110), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[5][37] ), .QN(n9109));
   SDFFARX1 \key_mem_reg[6][37]  (.D(n4782), .SI(n8982), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[6][37] ), .QN(n8981));
   SDFFARX1 \key_mem_reg[7][37]  (.D(n4783), .SI(n8854), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7366), .Q(\key_mem[7][37] ), .QN(n8853));
   SDFFARX1 \key_mem_reg[8][37]  (.D(n4784), .SI(n8726), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[8][37] ), .QN(n8725));
   SDFFARX1 \key_mem_reg[9][37]  (.D(n4785), .SI(n8598), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[9][37] ), .QN(n8597));
   SDFFARX1 \key_mem_reg[10][37]  (.D(n4786), .SI(n8470), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[10][37] ), .QN(n8469));
   SDFFARX1 \key_mem_reg[11][37]  (.D(n4787), .SI(n8342), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[11][37] ), .QN(n8341));
   SDFFARX1 \key_mem_reg[12][37]  (.D(n4788), .SI(n8214), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[12][37] ), .QN(n8213));
   SDFFARX1 \key_mem_reg[13][37]  (.D(n4789), .SI(n8087), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[13][37] ), .QN(n8086));
   SDFFARX1 \key_mem_reg[14][37]  (.D(n4790), .SI(n7959), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[14][37] ), .QN(n7958));
   SDFFARX1 \prev_key1_reg_reg[36]  (.D(n5437), .SI(n7720), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(prev_key1_reg[36]), .QN(n7719));
   SDFFARX1 \prev_key0_reg_reg[36]  (.D(n5564), .SI(n7832), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(prev_key0_reg[36]), .QN(n7831));
   SDFFARX1 \key_mem_reg[0][36]  (.D(n4791), .SI(n9750), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[0][36] ), .QN(n9749));
   SDFFARX1 \key_mem_reg[1][36]  (.D(n4792), .SI(n9622), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[1][36] ), .QN(n9621));
   SDFFARX1 \key_mem_reg[2][36]  (.D(n4793), .SI(n9494), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7365), .Q(\key_mem[2][36] ), .QN(n9493));
   SDFFARX1 \key_mem_reg[3][36]  (.D(n4794), .SI(n9366), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[3][36] ), .QN(n9365));
   SDFFARX1 \key_mem_reg[4][36]  (.D(n4795), .SI(n9238), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[4][36] ), .QN(n9237));
   SDFFARX1 \key_mem_reg[5][36]  (.D(n4796), .SI(n9111), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[5][36] ), .QN(n9110));
   SDFFARX1 \key_mem_reg[6][36]  (.D(n4797), .SI(n8983), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[6][36] ), .QN(n8982));
   SDFFARX1 \key_mem_reg[7][36]  (.D(n4798), .SI(n8855), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[7][36] ), .QN(n8854));
   SDFFARX1 \key_mem_reg[8][36]  (.D(n4799), .SI(n8727), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[8][36] ), .QN(n8726));
   SDFFARX1 \key_mem_reg[9][36]  (.D(n4800), .SI(n8599), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[9][36] ), .QN(n8598));
   SDFFARX1 \key_mem_reg[10][36]  (.D(n4801), .SI(n8471), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[10][36] ), .QN(n8470));
   SDFFARX1 \key_mem_reg[11][36]  (.D(n4802), .SI(n8343), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[11][36] ), .QN(n8342));
   SDFFARX1 \key_mem_reg[12][36]  (.D(n4803), .SI(n8215), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[12][36] ), .QN(n8214));
   SDFFARX1 \key_mem_reg[13][36]  (.D(n4804), .SI(n8088), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[13][36] ), .QN(n8087));
   SDFFARX1 \key_mem_reg[14][36]  (.D(n4805), .SI(n7960), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7364), .Q(\key_mem[14][36] ), .QN(n7959));
   SDFFARX1 \prev_key1_reg_reg[35]  (.D(n5438), .SI(n7721), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(prev_key1_reg[35]), .QN(n7720));
   SDFFARX1 \prev_key0_reg_reg[35]  (.D(n5565), .SI(n7833), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(prev_key0_reg[35]), .QN(n7832));
   SDFFARX1 \key_mem_reg[0][35]  (.D(n4806), .SI(n9751), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[0][35] ), .QN(n9750));
   SDFFARX1 \key_mem_reg[1][35]  (.D(n4807), .SI(n9623), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[1][35] ), .QN(n9622));
   SDFFARX1 \key_mem_reg[2][35]  (.D(n4808), .SI(n9495), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[2][35] ), .QN(n9494));
   SDFFARX1 \key_mem_reg[3][35]  (.D(n4809), .SI(n9367), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[3][35] ), .QN(n9366));
   SDFFARX1 \key_mem_reg[4][35]  (.D(n4810), .SI(n9239), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[4][35] ), .QN(n9238));
   SDFFARX1 \key_mem_reg[5][35]  (.D(n4811), .SI(n9112), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[5][35] ), .QN(n9111));
   SDFFARX1 \key_mem_reg[6][35]  (.D(n4812), .SI(n8984), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[6][35] ), .QN(n8983));
   SDFFARX1 \key_mem_reg[7][35]  (.D(n4813), .SI(n8856), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[7][35] ), .QN(n8855));
   SDFFARX1 \key_mem_reg[8][35]  (.D(n4814), .SI(n8728), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[8][35] ), .QN(n8727));
   SDFFARX1 \key_mem_reg[9][35]  (.D(n4815), .SI(n8600), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7363), .Q(\key_mem[9][35] ), .QN(n8599));
   SDFFARX1 \key_mem_reg[10][35]  (.D(n4816), .SI(n8472), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[10][35] ), .QN(n8471));
   SDFFARX1 \key_mem_reg[11][35]  (.D(n4817), .SI(n8344), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[11][35] ), .QN(n8343));
   SDFFARX1 \key_mem_reg[12][35]  (.D(n4818), .SI(n8216), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[12][35] ), .QN(n8215));
   SDFFARX1 \key_mem_reg[13][35]  (.D(n4819), .SI(n8089), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[13][35] ), .QN(n8088));
   SDFFARX1 \key_mem_reg[14][35]  (.D(n4820), .SI(n7961), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[14][35] ), .QN(n7960));
   SDFFARX1 \prev_key1_reg_reg[34]  (.D(n5439), .SI(n7722), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(prev_key1_reg[34]), .QN(n7721));
   SDFFARX1 \prev_key0_reg_reg[34]  (.D(n5566), .SI(n7834), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(prev_key0_reg[34]), .QN(n7833));
   SDFFARX1 \key_mem_reg[0][34]  (.D(n4821), .SI(n9752), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[0][34] ), .QN(n9751));
   SDFFARX1 \key_mem_reg[1][34]  (.D(n4822), .SI(n9624), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[1][34] ), .QN(n9623));
   SDFFARX1 \key_mem_reg[2][34]  (.D(n4823), .SI(n9496), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[2][34] ), .QN(n9495));
   SDFFARX1 \key_mem_reg[3][34]  (.D(n4824), .SI(n9368), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[3][34] ), .QN(n9367));
   SDFFARX1 \key_mem_reg[4][34]  (.D(n4825), .SI(n9240), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7362), .Q(\key_mem[4][34] ), .QN(n9239));
   SDFFARX1 \key_mem_reg[5][34]  (.D(n4826), .SI(n9113), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[5][34] ), .QN(n9112));
   SDFFARX1 \key_mem_reg[6][34]  (.D(n4827), .SI(n8985), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[6][34] ), .QN(n8984));
   SDFFARX1 \key_mem_reg[7][34]  (.D(n4828), .SI(n8857), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[7][34] ), .QN(n8856));
   SDFFARX1 \key_mem_reg[8][34]  (.D(n4829), .SI(n8729), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[8][34] ), .QN(n8728));
   SDFFARX1 \key_mem_reg[9][34]  (.D(n4830), .SI(n8601), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[9][34] ), .QN(n8600));
   SDFFARX1 \key_mem_reg[10][34]  (.D(n4831), .SI(n8473), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[10][34] ), .QN(n8472));
   SDFFARX1 \key_mem_reg[11][34]  (.D(n4832), .SI(n8345), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[11][34] ), .QN(n8344));
   SDFFARX1 \key_mem_reg[12][34]  (.D(n4833), .SI(n8217), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[12][34] ), .QN(n8216));
   SDFFARX1 \key_mem_reg[13][34]  (.D(n4834), .SI(n8090), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[13][34] ), .QN(n8089));
   SDFFARX1 \key_mem_reg[14][34]  (.D(n4835), .SI(n7962), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(\key_mem[14][34] ), .QN(n7961));
   SDFFARX1 \prev_key1_reg_reg[33]  (.D(n5440), .SI(n7723), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(prev_key1_reg[33]), .QN(n7722));
   SDFFARX1 \prev_key0_reg_reg[33]  (.D(n5567), .SI(n7835), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7361), .Q(prev_key0_reg[33]), .QN(n7834));
   SDFFARX1 \key_mem_reg[0][33]  (.D(n4836), .SI(n9753), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[0][33] ), .QN(n9752));
   SDFFARX1 \key_mem_reg[1][33]  (.D(n4837), .SI(n9625), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[1][33] ), .QN(n9624));
   SDFFARX1 \key_mem_reg[2][33]  (.D(n4838), .SI(n9497), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[2][33] ), .QN(n9496));
   SDFFARX1 \key_mem_reg[3][33]  (.D(n4839), .SI(n9369), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[3][33] ), .QN(n9368));
   SDFFARX1 \key_mem_reg[4][33]  (.D(n4840), .SI(n9241), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[4][33] ), .QN(n9240));
   SDFFARX1 \key_mem_reg[5][33]  (.D(n4841), .SI(n9114), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[5][33] ), .QN(n9113));
   SDFFARX1 \key_mem_reg[6][33]  (.D(n4842), .SI(n8986), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[6][33] ), .QN(n8985));
   SDFFARX1 \key_mem_reg[7][33]  (.D(n4843), .SI(n8858), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[7][33] ), .QN(n8857));
   SDFFARX1 \key_mem_reg[8][33]  (.D(n4844), .SI(n8730), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[8][33] ), .QN(n8729));
   SDFFARX1 \key_mem_reg[9][33]  (.D(n4845), .SI(n8602), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[9][33] ), .QN(n8601));
   SDFFARX1 \key_mem_reg[10][33]  (.D(n4846), .SI(n8474), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[10][33] ), .QN(n8473));
   SDFFARX1 \key_mem_reg[11][33]  (.D(n4847), .SI(n8346), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7360), .Q(\key_mem[11][33] ), .QN(n8345));
   SDFFARX1 \key_mem_reg[12][33]  (.D(n4848), .SI(n8218), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[12][33] ), .QN(n8217));
   SDFFARX1 \key_mem_reg[13][33]  (.D(n4849), .SI(n8091), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[13][33] ), .QN(n8090));
   SDFFARX1 \key_mem_reg[14][33]  (.D(n4850), .SI(n7963), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[14][33] ), .QN(n7962));
   SDFFARX1 \prev_key1_reg_reg[32]  (.D(n5441), .SI(n7724), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(prev_key1_reg[32]), .QN(n7723));
   SDFFARX1 \prev_key0_reg_reg[32]  (.D(n5568), .SI(n7836), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(prev_key0_reg[32]), .QN(n7835));
   SDFFARX1 \key_mem_reg[0][32]  (.D(n4851), .SI(n9754), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[0][32] ), .QN(n9753));
   SDFFARX1 \key_mem_reg[1][32]  (.D(n4852), .SI(n9626), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[1][32] ), .QN(n9625));
   SDFFARX1 \key_mem_reg[2][32]  (.D(n4853), .SI(n9498), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[2][32] ), .QN(n9497));
   SDFFARX1 \key_mem_reg[3][32]  (.D(n4854), .SI(n9370), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[3][32] ), .QN(n9369));
   SDFFARX1 \key_mem_reg[4][32]  (.D(n4855), .SI(n9242), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[4][32] ), .QN(n9241));
   SDFFARX1 \key_mem_reg[5][32]  (.D(n4856), .SI(n9115), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[5][32] ), .QN(n9114));
   SDFFARX1 \key_mem_reg[6][32]  (.D(n4857), .SI(n8987), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7359), .Q(\key_mem[6][32] ), .QN(n8986));
   SDFFARX1 \key_mem_reg[7][32]  (.D(n4858), .SI(n8859), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[7][32] ), .QN(n8858));
   SDFFARX1 \key_mem_reg[8][32]  (.D(n4859), .SI(n8731), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[8][32] ), .QN(n8730));
   SDFFARX1 \key_mem_reg[9][32]  (.D(n4860), .SI(n8603), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[9][32] ), .QN(n8602));
   SDFFARX1 \key_mem_reg[10][32]  (.D(n4861), .SI(n8475), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[10][32] ), .QN(n8474));
   SDFFARX1 \key_mem_reg[11][32]  (.D(n4862), .SI(n8347), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[11][32] ), .QN(n8346));
   SDFFARX1 \key_mem_reg[12][32]  (.D(n4863), .SI(n8219), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[12][32] ), .QN(n8218));
   SDFFARX1 \key_mem_reg[13][32]  (.D(n4864), .SI(n8092), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[13][32] ), .QN(n8091));
   SDFFARX1 \key_mem_reg[14][32]  (.D(n4865), .SI(n7964), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[14][32] ), .QN(n7963));
   SDFFARX1 \prev_key1_reg_reg[31]  (.D(n5442), .SI(n7725), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(sboxw[31]), .QN(n7724));
   SDFFARX1 \prev_key0_reg_reg[31]  (.D(n5569), .SI(n7837), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(prev_key0_reg[31]), .QN(n7836));
   SDFFARX1 \key_mem_reg[0][31]  (.D(n4866), .SI(n9755), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[0][31] ), .QN(n9754));
   SDFFARX1 \key_mem_reg[1][31]  (.D(n4867), .SI(n9627), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7358), .Q(\key_mem[1][31] ), .QN(n9626));
   SDFFARX1 \key_mem_reg[2][31]  (.D(n4868), .SI(n9499), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[2][31] ), .QN(n9498));
   SDFFARX1 \key_mem_reg[3][31]  (.D(n4869), .SI(n9371), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[3][31] ), .QN(n9370));
   SDFFARX1 \key_mem_reg[4][31]  (.D(n4870), .SI(n9243), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[4][31] ), .QN(n9242));
   SDFFARX1 \key_mem_reg[5][31]  (.D(n4871), .SI(n9116), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[5][31] ), .QN(n9115));
   SDFFARX1 \key_mem_reg[6][31]  (.D(n4872), .SI(n8988), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[6][31] ), .QN(n8987));
   SDFFARX1 \key_mem_reg[7][31]  (.D(n4873), .SI(n8860), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[7][31] ), .QN(n8859));
   SDFFARX1 \key_mem_reg[8][31]  (.D(n4874), .SI(n8732), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[8][31] ), .QN(n8731));
   SDFFARX1 \key_mem_reg[9][31]  (.D(n4875), .SI(n8604), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[9][31] ), .QN(n8603));
   SDFFARX1 \key_mem_reg[10][31]  (.D(n4876), .SI(n8476), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[10][31] ), .QN(n8475));
   SDFFARX1 \key_mem_reg[11][31]  (.D(n4877), .SI(n8348), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[11][31] ), .QN(n8347));
   SDFFARX1 \key_mem_reg[12][31]  (.D(n4878), .SI(n8220), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[12][31] ), .QN(n8219));
   SDFFARX1 \key_mem_reg[13][31]  (.D(n4879), .SI(n8093), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7357), .Q(\key_mem[13][31] ), .QN(n8092));
   SDFFARX1 \key_mem_reg[14][31]  (.D(n4880), .SI(n7965), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[14][31] ), .QN(n7964));
   SDFFARX1 \prev_key1_reg_reg[30]  (.D(n5443), .SI(n7726), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(sboxw[30]), .QN(n7725));
   SDFFARX1 \prev_key0_reg_reg[30]  (.D(n5570), .SI(n7838), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(prev_key0_reg[30]), .QN(n7837));
   SDFFARX1 \key_mem_reg[0][30]  (.D(n4881), .SI(n9756), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[0][30] ), .QN(n9755));
   SDFFARX1 \key_mem_reg[1][30]  (.D(n4882), .SI(n9628), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[1][30] ), .QN(n9627));
   SDFFARX1 \key_mem_reg[2][30]  (.D(n4883), .SI(n9500), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[2][30] ), .QN(n9499));
   SDFFARX1 \key_mem_reg[3][30]  (.D(n4884), .SI(n9372), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[3][30] ), .QN(n9371));
   SDFFARX1 \key_mem_reg[4][30]  (.D(n4885), .SI(n9244), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[4][30] ), .QN(n9243));
   SDFFARX1 \key_mem_reg[5][30]  (.D(n4886), .SI(n9117), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[5][30] ), .QN(n9116));
   SDFFARX1 \key_mem_reg[6][30]  (.D(n4887), .SI(n8989), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[6][30] ), .QN(n8988));
   SDFFARX1 \key_mem_reg[7][30]  (.D(n4888), .SI(n8861), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[7][30] ), .QN(n8860));
   SDFFARX1 \key_mem_reg[8][30]  (.D(n4889), .SI(n8733), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7356), .Q(\key_mem[8][30] ), .QN(n8732));
   SDFFARX1 \key_mem_reg[9][30]  (.D(n4890), .SI(n8605), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[9][30] ), .QN(n8604));
   SDFFARX1 \key_mem_reg[10][30]  (.D(n4891), .SI(n8477), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[10][30] ), .QN(n8476));
   SDFFARX1 \key_mem_reg[11][30]  (.D(n4892), .SI(n8349), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[11][30] ), .QN(n8348));
   SDFFARX1 \key_mem_reg[12][30]  (.D(n4893), .SI(n8221), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[12][30] ), .QN(n8220));
   SDFFARX1 \key_mem_reg[13][30]  (.D(n4894), .SI(n8094), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[13][30] ), .QN(n8093));
   SDFFARX1 \key_mem_reg[14][30]  (.D(n4895), .SI(n7966), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[14][30] ), .QN(n7965));
   SDFFARX1 \prev_key1_reg_reg[29]  (.D(n5444), .SI(n7727), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(sboxw[29]), .QN(n7726));
   SDFFARX1 \prev_key0_reg_reg[29]  (.D(n5571), .SI(n7839), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(prev_key0_reg[29]), .QN(n7838));
   SDFFARX1 \key_mem_reg[0][29]  (.D(n4896), .SI(n9757), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[0][29] ), .QN(n9756));
   SDFFARX1 \key_mem_reg[1][29]  (.D(n4897), .SI(n9629), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[1][29] ), .QN(n9628));
   SDFFARX1 \key_mem_reg[2][29]  (.D(n4898), .SI(n9501), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[2][29] ), .QN(n9500));
   SDFFARX1 \key_mem_reg[3][29]  (.D(n4899), .SI(n9373), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7355), .Q(\key_mem[3][29] ), .QN(n9372));
   SDFFARX1 \key_mem_reg[4][29]  (.D(n4900), .SI(n9245), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[4][29] ), .QN(n9244));
   SDFFARX1 \key_mem_reg[5][29]  (.D(n4901), .SI(n9118), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[5][29] ), .QN(n9117));
   SDFFARX1 \key_mem_reg[6][29]  (.D(n4902), .SI(n8990), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[6][29] ), .QN(n8989));
   SDFFARX1 \key_mem_reg[7][29]  (.D(n4903), .SI(n8862), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[7][29] ), .QN(n8861));
   SDFFARX1 \key_mem_reg[8][29]  (.D(n4904), .SI(n8734), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[8][29] ), .QN(n8733));
   SDFFARX1 \key_mem_reg[9][29]  (.D(n4905), .SI(n8606), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[9][29] ), .QN(n8605));
   SDFFARX1 \key_mem_reg[10][29]  (.D(n4906), .SI(n8478), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[10][29] ), .QN(n8477));
   SDFFARX1 \key_mem_reg[11][29]  (.D(n4907), .SI(n8350), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[11][29] ), .QN(n8349));
   SDFFARX1 \key_mem_reg[12][29]  (.D(n4908), .SI(n8222), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[12][29] ), .QN(n8221));
   SDFFARX1 \key_mem_reg[13][29]  (.D(n4909), .SI(n8095), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[13][29] ), .QN(n8094));
   SDFFARX1 \key_mem_reg[14][29]  (.D(n4910), .SI(n7967), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(\key_mem[14][29] ), .QN(n7966));
   SDFFARX1 \prev_key1_reg_reg[28]  (.D(n5445), .SI(n7728), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7354), .Q(sboxw[28]), .QN(n7727));
   SDFFARX1 \prev_key0_reg_reg[28]  (.D(n5572), .SI(n7840), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(prev_key0_reg[28]), .QN(n7839));
   SDFFARX1 \key_mem_reg[0][28]  (.D(n4911), .SI(n9758), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[0][28] ), .QN(n9757));
   SDFFARX1 \key_mem_reg[1][28]  (.D(n4912), .SI(n9630), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[1][28] ), .QN(n9629));
   SDFFARX1 \key_mem_reg[2][28]  (.D(n4913), .SI(n9502), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[2][28] ), .QN(n9501));
   SDFFARX1 \key_mem_reg[3][28]  (.D(n4914), .SI(n9374), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[3][28] ), .QN(n9373));
   SDFFARX1 \key_mem_reg[4][28]  (.D(n4915), .SI(n9246), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[4][28] ), .QN(n9245));
   SDFFARX1 \key_mem_reg[5][28]  (.D(n4916), .SI(n9119), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[5][28] ), .QN(n9118));
   SDFFARX1 \key_mem_reg[6][28]  (.D(n4917), .SI(n8991), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[6][28] ), .QN(n8990));
   SDFFARX1 \key_mem_reg[7][28]  (.D(n4918), .SI(n8863), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[7][28] ), .QN(n8862));
   SDFFARX1 \key_mem_reg[8][28]  (.D(n4919), .SI(n8735), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[8][28] ), .QN(n8734));
   SDFFARX1 \key_mem_reg[9][28]  (.D(n4920), .SI(n8607), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[9][28] ), .QN(n8606));
   SDFFARX1 \key_mem_reg[10][28]  (.D(n4921), .SI(n8479), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7353), .Q(\key_mem[10][28] ), .QN(n8478));
   SDFFARX1 \key_mem_reg[11][28]  (.D(n4922), .SI(n8351), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[11][28] ), .QN(n8350));
   SDFFARX1 \key_mem_reg[12][28]  (.D(n4923), .SI(n8223), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[12][28] ), .QN(n8222));
   SDFFARX1 \key_mem_reg[13][28]  (.D(n4924), .SI(n8096), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[13][28] ), .QN(n8095));
   SDFFARX1 \key_mem_reg[14][28]  (.D(n4925), .SI(n7968), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[14][28] ), .QN(n7967));
   SDFFARX1 \prev_key1_reg_reg[27]  (.D(n5446), .SI(n7729), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(sboxw[27]), .QN(n7728));
   SDFFARX1 \prev_key0_reg_reg[27]  (.D(n5573), .SI(n7841), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(prev_key0_reg[27]), .QN(n7840));
   SDFFARX1 \key_mem_reg[0][27]  (.D(n4926), .SI(n9759), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[0][27] ), .QN(n9758));
   SDFFARX1 \key_mem_reg[1][27]  (.D(n4927), .SI(n9631), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[1][27] ), .QN(n9630));
   SDFFARX1 \key_mem_reg[2][27]  (.D(n4928), .SI(n9503), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[2][27] ), .QN(n9502));
   SDFFARX1 \key_mem_reg[3][27]  (.D(n4929), .SI(n9375), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[3][27] ), .QN(n9374));
   SDFFARX1 \key_mem_reg[4][27]  (.D(n4930), .SI(n9247), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[4][27] ), .QN(n9246));
   SDFFARX1 \key_mem_reg[5][27]  (.D(n4931), .SI(n9120), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7352), .Q(\key_mem[5][27] ), .QN(n9119));
   SDFFARX1 \key_mem_reg[6][27]  (.D(n4932), .SI(n8992), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[6][27] ), .QN(n8991));
   SDFFARX1 \key_mem_reg[7][27]  (.D(n4933), .SI(n8864), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[7][27] ), .QN(n8863));
   SDFFARX1 \key_mem_reg[8][27]  (.D(n4934), .SI(n8736), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[8][27] ), .QN(n8735));
   SDFFARX1 \key_mem_reg[9][27]  (.D(n4935), .SI(n8608), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[9][27] ), .QN(n8607));
   SDFFARX1 \key_mem_reg[10][27]  (.D(n4936), .SI(n8480), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[10][27] ), .QN(n8479));
   SDFFARX1 \key_mem_reg[11][27]  (.D(n4937), .SI(n8352), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[11][27] ), .QN(n8351));
   SDFFARX1 \key_mem_reg[12][27]  (.D(n4938), .SI(n8224), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[12][27] ), .QN(n8223));
   SDFFARX1 \key_mem_reg[13][27]  (.D(n4939), .SI(n8097), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[13][27] ), .QN(n8096));
   SDFFARX1 \key_mem_reg[14][27]  (.D(n4940), .SI(n7969), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[14][27] ), .QN(n7968));
   SDFFARX1 \prev_key1_reg_reg[26]  (.D(n5447), .SI(n7730), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(sboxw[26]), .QN(n7729));
   SDFFARX1 \prev_key0_reg_reg[26]  (.D(n5574), .SI(n7842), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(prev_key0_reg[26]), .QN(n7841));
   SDFFARX1 \key_mem_reg[0][26]  (.D(n4941), .SI(n9760), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7351), .Q(\key_mem[0][26] ), .QN(n9759));
   SDFFARX1 \key_mem_reg[1][26]  (.D(n4942), .SI(n9632), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[1][26] ), .QN(n9631));
   SDFFARX1 \key_mem_reg[2][26]  (.D(n4943), .SI(n9504), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[2][26] ), .QN(n9503));
   SDFFARX1 \key_mem_reg[3][26]  (.D(n4944), .SI(n9376), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[3][26] ), .QN(n9375));
   SDFFARX1 \key_mem_reg[4][26]  (.D(n4945), .SI(n9248), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[4][26] ), .QN(n9247));
   SDFFARX1 \key_mem_reg[5][26]  (.D(n4946), .SI(n9121), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[5][26] ), .QN(n9120));
   SDFFARX1 \key_mem_reg[6][26]  (.D(n4947), .SI(n8993), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[6][26] ), .QN(n8992));
   SDFFARX1 \key_mem_reg[7][26]  (.D(n4948), .SI(n8865), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[7][26] ), .QN(n8864));
   SDFFARX1 \key_mem_reg[8][26]  (.D(n4949), .SI(n8737), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[8][26] ), .QN(n8736));
   SDFFARX1 \key_mem_reg[9][26]  (.D(n4950), .SI(n8609), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[9][26] ), .QN(n8608));
   SDFFARX1 \key_mem_reg[10][26]  (.D(n4951), .SI(n8481), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[10][26] ), .QN(n8480));
   SDFFARX1 \key_mem_reg[11][26]  (.D(n4952), .SI(n8353), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[11][26] ), .QN(n8352));
   SDFFARX1 \key_mem_reg[12][26]  (.D(n4953), .SI(n8225), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7350), .Q(\key_mem[12][26] ), .QN(n8224));
   SDFFARX1 \key_mem_reg[13][26]  (.D(n4954), .SI(n8098), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[13][26] ), .QN(n8097));
   SDFFARX1 \key_mem_reg[14][26]  (.D(n4955), .SI(n7970), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[14][26] ), .QN(n7969));
   SDFFARX1 \prev_key1_reg_reg[25]  (.D(n5448), .SI(n7731), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(sboxw[25]), .QN(n7730));
   SDFFARX1 \prev_key0_reg_reg[25]  (.D(n5575), .SI(n7843), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(prev_key0_reg[25]), .QN(n7842));
   SDFFARX1 \key_mem_reg[0][25]  (.D(n4956), .SI(n9761), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[0][25] ), .QN(n9760));
   SDFFARX1 \key_mem_reg[1][25]  (.D(n4957), .SI(n9633), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[1][25] ), .QN(n9632));
   SDFFARX1 \key_mem_reg[2][25]  (.D(n4958), .SI(n9505), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[2][25] ), .QN(n9504));
   SDFFARX1 \key_mem_reg[3][25]  (.D(n4959), .SI(n9377), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[3][25] ), .QN(n9376));
   SDFFARX1 \key_mem_reg[4][25]  (.D(n4960), .SI(n9249), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[4][25] ), .QN(n9248));
   SDFFARX1 \key_mem_reg[5][25]  (.D(n4961), .SI(n9122), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[5][25] ), .QN(n9121));
   SDFFARX1 \key_mem_reg[6][25]  (.D(n4962), .SI(n8994), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[6][25] ), .QN(n8993));
   SDFFARX1 \key_mem_reg[7][25]  (.D(n4963), .SI(n8866), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7349), .Q(\key_mem[7][25] ), .QN(n8865));
   SDFFARX1 \key_mem_reg[8][25]  (.D(n4964), .SI(n8738), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[8][25] ), .QN(n8737));
   SDFFARX1 \key_mem_reg[9][25]  (.D(n4965), .SI(n8610), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[9][25] ), .QN(n8609));
   SDFFARX1 \key_mem_reg[10][25]  (.D(n4966), .SI(n8482), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[10][25] ), .QN(n8481));
   SDFFARX1 \key_mem_reg[11][25]  (.D(n4967), .SI(n8354), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[11][25] ), .QN(n8353));
   SDFFARX1 \key_mem_reg[12][25]  (.D(n4968), .SI(n8226), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[12][25] ), .QN(n8225));
   SDFFARX1 \key_mem_reg[13][25]  (.D(n4969), .SI(n8099), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[13][25] ), .QN(n8098));
   SDFFARX1 \key_mem_reg[14][25]  (.D(n4970), .SI(n7971), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[14][25] ), .QN(n7970));
   SDFFARX1 \prev_key1_reg_reg[24]  (.D(n5449), .SI(n7732), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(sboxw[24]), .QN(n7731));
   SDFFARX1 \prev_key0_reg_reg[24]  (.D(n5576), .SI(n7844), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(prev_key0_reg[24]), .QN(n7843));
   SDFFARX1 \key_mem_reg[0][24]  (.D(n4971), .SI(n9762), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[0][24] ), .QN(n9761));
   SDFFARX1 \key_mem_reg[1][24]  (.D(n4972), .SI(n9634), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[1][24] ), .QN(n9633));
   SDFFARX1 \key_mem_reg[2][24]  (.D(n4973), .SI(n9506), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7348), .Q(\key_mem[2][24] ), .QN(n9505));
   SDFFARX1 \key_mem_reg[3][24]  (.D(n4974), .SI(n9378), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[3][24] ), .QN(n9377));
   SDFFARX1 \key_mem_reg[4][24]  (.D(n4975), .SI(n9250), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[4][24] ), .QN(n9249));
   SDFFARX1 \key_mem_reg[5][24]  (.D(n4976), .SI(n9123), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[5][24] ), .QN(n9122));
   SDFFARX1 \key_mem_reg[6][24]  (.D(n4977), .SI(n8995), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[6][24] ), .QN(n8994));
   SDFFARX1 \key_mem_reg[7][24]  (.D(n4978), .SI(n8867), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[7][24] ), .QN(n8866));
   SDFFARX1 \key_mem_reg[8][24]  (.D(n4979), .SI(n8739), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[8][24] ), .QN(n8738));
   SDFFARX1 \key_mem_reg[9][24]  (.D(n4980), .SI(n8611), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[9][24] ), .QN(n8610));
   SDFFARX1 \key_mem_reg[10][24]  (.D(n4981), .SI(n8483), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[10][24] ), .QN(n8482));
   SDFFARX1 \key_mem_reg[11][24]  (.D(n4982), .SI(n8355), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[11][24] ), .QN(n8354));
   SDFFARX1 \key_mem_reg[12][24]  (.D(n4983), .SI(n8227), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[12][24] ), .QN(n8226));
   SDFFARX1 \key_mem_reg[13][24]  (.D(n4984), .SI(n8100), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[13][24] ), .QN(n8099));
   SDFFARX1 \key_mem_reg[14][24]  (.D(n4985), .SI(n7972), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7347), .Q(\key_mem[14][24] ), .QN(n7971));
   SDFFARX1 \prev_key1_reg_reg[23]  (.D(n5450), .SI(n7733), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(sboxw[23]), .QN(n7732));
   SDFFARX1 \prev_key0_reg_reg[23]  (.D(n5577), .SI(n7845), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(prev_key0_reg[23]), .QN(n7844));
   SDFFARX1 \key_mem_reg[0][23]  (.D(n4986), .SI(n9763), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(\key_mem[0][23] ), .QN(n9762));
   SDFFARX1 \key_mem_reg[1][23]  (.D(n4987), .SI(n9635), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(\key_mem[1][23] ), .QN(n9634));
   SDFFARX1 \key_mem_reg[2][23]  (.D(n4988), .SI(n9507), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(\key_mem[2][23] ), .QN(n9506));
   SDFFARX1 \key_mem_reg[3][23]  (.D(n4989), .SI(n9379), .SE(test_se_buf_net5), .CLK(
          clk_buf_net5), .RSTB(n7346), .Q(\key_mem[3][23] ), .QN(n9378));
   SDFFARX1 \key_mem_reg[4][23]  (.D(n4990), .SI(n9251), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[4][23] ), .QN(n9250));
   SDFFARX1 \key_mem_reg[5][23]  (.D(n4991), .SI(n9124), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[5][23] ), .QN(n9123));
   SDFFARX1 \key_mem_reg[6][23]  (.D(n4992), .SI(n8996), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[6][23] ), .QN(n8995));
   SDFFARX1 \key_mem_reg[7][23]  (.D(n4993), .SI(n8868), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[7][23] ), .QN(n8867));
   SDFFARX1 \key_mem_reg[8][23]  (.D(n4994), .SI(n8740), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[8][23] ), .QN(n8739));
   SDFFARX1 \key_mem_reg[9][23]  (.D(n4995), .SI(n8612), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7346), .Q(\key_mem[9][23] ), .QN(n8611));
   SDFFARX1 \key_mem_reg[10][23]  (.D(n4996), .SI(n8484), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[10][23] ), .QN(n8483));
   SDFFARX1 \key_mem_reg[11][23]  (.D(n4997), .SI(n8356), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[11][23] ), .QN(n8355));
   SDFFARX1 \key_mem_reg[12][23]  (.D(n4998), .SI(n8228), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[12][23] ), .QN(n8227));
   SDFFARX1 \key_mem_reg[13][23]  (.D(n4999), .SI(n8101), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[13][23] ), .QN(n8100));
   SDFFARX1 \key_mem_reg[14][23]  (.D(n5000), .SI(n7973), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[14][23] ), .QN(n7972));
   SDFFARX1 \prev_key1_reg_reg[22]  (.D(n5451), .SI(n7734), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(sboxw[22]), .QN(n7733));
   SDFFARX1 \prev_key0_reg_reg[22]  (.D(n5578), .SI(n7846), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(prev_key0_reg[22]), .QN(n7845));
   SDFFARX1 \key_mem_reg[0][22]  (.D(n5001), .SI(n9764), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[0][22] ), .QN(n9763));
   SDFFARX1 \key_mem_reg[1][22]  (.D(n5002), .SI(n9636), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[1][22] ), .QN(n9635));
   SDFFARX1 \key_mem_reg[2][22]  (.D(n5003), .SI(n9508), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[2][22] ), .QN(n9507));
   SDFFARX1 \key_mem_reg[3][22]  (.D(n5004), .SI(n9380), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[3][22] ), .QN(n9379));
   SDFFARX1 \key_mem_reg[4][22]  (.D(n5005), .SI(n9252), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7345), .Q(\key_mem[4][22] ), .QN(n9251));
   SDFFARX1 \key_mem_reg[5][22]  (.D(n5006), .SI(n9125), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[5][22] ), .QN(n9124));
   SDFFARX1 \key_mem_reg[6][22]  (.D(n5007), .SI(n8997), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[6][22] ), .QN(n8996));
   SDFFARX1 \key_mem_reg[7][22]  (.D(n5008), .SI(n8869), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[7][22] ), .QN(n8868));
   SDFFARX1 \key_mem_reg[8][22]  (.D(n5009), .SI(n8741), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[8][22] ), .QN(n8740));
   SDFFARX1 \key_mem_reg[9][22]  (.D(n5010), .SI(n8613), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[9][22] ), .QN(n8612));
   SDFFARX1 \key_mem_reg[10][22]  (.D(n5011), .SI(n8485), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[10][22] ), .QN(n8484));
   SDFFARX1 \key_mem_reg[11][22]  (.D(n5012), .SI(n8357), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[11][22] ), .QN(n8356));
   SDFFARX1 \key_mem_reg[12][22]  (.D(n5013), .SI(n8229), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[12][22] ), .QN(n8228));
   SDFFARX1 \key_mem_reg[13][22]  (.D(n5014), .SI(n8102), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[13][22] ), .QN(n8101));
   SDFFARX1 \key_mem_reg[14][22]  (.D(n5015), .SI(n7974), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(\key_mem[14][22] ), .QN(n7973));
   SDFFARX1 \prev_key1_reg_reg[21]  (.D(n5452), .SI(n7735), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(sboxw[21]), .QN(n7734));
   SDFFARX1 \prev_key0_reg_reg[21]  (.D(n5579), .SI(n7847), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7344), .Q(prev_key0_reg[21]), .QN(n7846));
   SDFFARX1 \key_mem_reg[0][21]  (.D(n5016), .SI(n9765), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[0][21] ), .QN(n9764));
   SDFFARX1 \key_mem_reg[1][21]  (.D(n5017), .SI(n9637), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[1][21] ), .QN(n9636));
   SDFFARX1 \key_mem_reg[2][21]  (.D(n5018), .SI(n9509), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[2][21] ), .QN(n9508));
   SDFFARX1 \key_mem_reg[3][21]  (.D(n5019), .SI(n9381), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[3][21] ), .QN(n9380));
   SDFFARX1 \key_mem_reg[4][21]  (.D(n5020), .SI(n9253), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[4][21] ), .QN(n9252));
   SDFFARX1 \key_mem_reg[5][21]  (.D(n5021), .SI(n9126), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[5][21] ), .QN(n9125));
   SDFFARX1 \key_mem_reg[6][21]  (.D(n5022), .SI(n8998), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[6][21] ), .QN(n8997));
   SDFFARX1 \key_mem_reg[7][21]  (.D(n5023), .SI(n8870), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[7][21] ), .QN(n8869));
   SDFFARX1 \key_mem_reg[8][21]  (.D(n5024), .SI(n8742), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[8][21] ), .QN(n8741));
   SDFFARX1 \key_mem_reg[9][21]  (.D(n5025), .SI(n8614), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[9][21] ), .QN(n8613));
   SDFFARX1 \key_mem_reg[10][21]  (.D(n5026), .SI(n8486), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[10][21] ), .QN(n8485));
   SDFFARX1 \key_mem_reg[11][21]  (.D(n5027), .SI(n8358), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7343), .Q(\key_mem[11][21] ), .QN(n8357));
   SDFFARX1 \key_mem_reg[12][21]  (.D(n5028), .SI(n8230), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[12][21] ), .QN(n8229));
   SDFFARX1 \key_mem_reg[13][21]  (.D(n5029), .SI(n8103), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[13][21] ), .QN(n8102));
   SDFFARX1 \key_mem_reg[14][21]  (.D(n5030), .SI(n7975), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[14][21] ), .QN(n7974));
   SDFFARX1 \prev_key1_reg_reg[20]  (.D(n5453), .SI(n7736), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(sboxw[20]), .QN(n7735));
   SDFFARX1 \prev_key0_reg_reg[20]  (.D(n5580), .SI(n7848), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(prev_key0_reg[20]), .QN(n7847));
   SDFFARX1 \key_mem_reg[0][20]  (.D(n5031), .SI(n9766), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[0][20] ), .QN(n9765));
   SDFFARX1 \key_mem_reg[1][20]  (.D(n5032), .SI(n9638), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[1][20] ), .QN(n9637));
   SDFFARX1 \key_mem_reg[2][20]  (.D(n5033), .SI(n9510), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[2][20] ), .QN(n9509));
   SDFFARX1 \key_mem_reg[3][20]  (.D(n5034), .SI(n9382), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[3][20] ), .QN(n9381));
   SDFFARX1 \key_mem_reg[4][20]  (.D(n5035), .SI(n9254), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[4][20] ), .QN(n9253));
   SDFFARX1 \key_mem_reg[5][20]  (.D(n5036), .SI(n9127), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[5][20] ), .QN(n9126));
   SDFFARX1 \key_mem_reg[6][20]  (.D(n5037), .SI(n8999), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7342), .Q(\key_mem[6][20] ), .QN(n8998));
   SDFFARX1 \key_mem_reg[7][20]  (.D(n5038), .SI(n8871), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[7][20] ), .QN(n8870));
   SDFFARX1 \key_mem_reg[8][20]  (.D(n5039), .SI(n8743), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[8][20] ), .QN(n8742));
   SDFFARX1 \key_mem_reg[9][20]  (.D(n5040), .SI(n8615), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[9][20] ), .QN(n8614));
   SDFFARX1 \key_mem_reg[10][20]  (.D(n5041), .SI(n8487), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[10][20] ), .QN(n8486));
   SDFFARX1 \key_mem_reg[11][20]  (.D(n5042), .SI(n8359), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[11][20] ), .QN(n8358));
   SDFFARX1 \key_mem_reg[12][20]  (.D(n5043), .SI(n8231), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[12][20] ), .QN(n8230));
   SDFFARX1 \key_mem_reg[13][20]  (.D(n5044), .SI(n8104), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[13][20] ), .QN(n8103));
   SDFFARX1 \key_mem_reg[14][20]  (.D(n5045), .SI(n7976), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[14][20] ), .QN(n7975));
   SDFFARX1 \prev_key1_reg_reg[19]  (.D(n5454), .SI(n7737), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(sboxw[19]), .QN(n7736));
   SDFFARX1 \prev_key0_reg_reg[19]  (.D(n5581), .SI(n7849), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(prev_key0_reg[19]), .QN(n7848));
   SDFFARX1 \key_mem_reg[0][19]  (.D(n5046), .SI(n9767), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[0][19] ), .QN(n9766));
   SDFFARX1 \key_mem_reg[1][19]  (.D(n5047), .SI(n9639), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7341), .Q(\key_mem[1][19] ), .QN(n9638));
   SDFFARX1 \key_mem_reg[2][19]  (.D(n5048), .SI(n9511), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[2][19] ), .QN(n9510));
   SDFFARX1 \key_mem_reg[3][19]  (.D(n5049), .SI(n9383), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[3][19] ), .QN(n9382));
   SDFFARX1 \key_mem_reg[4][19]  (.D(n5050), .SI(n9255), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[4][19] ), .QN(n9254));
   SDFFARX1 \key_mem_reg[5][19]  (.D(n5051), .SI(n9128), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[5][19] ), .QN(n9127));
   SDFFARX1 \key_mem_reg[6][19]  (.D(n5052), .SI(n9000), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[6][19] ), .QN(n8999));
   SDFFARX1 \key_mem_reg[7][19]  (.D(n5053), .SI(n8872), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[7][19] ), .QN(n8871));
   SDFFARX1 \key_mem_reg[8][19]  (.D(n5054), .SI(n8744), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[8][19] ), .QN(n8743));
   SDFFARX1 \key_mem_reg[9][19]  (.D(n5055), .SI(n8616), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[9][19] ), .QN(n8615));
   SDFFARX1 \key_mem_reg[10][19]  (.D(n5056), .SI(n8488), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[10][19] ), .QN(n8487));
   SDFFARX1 \key_mem_reg[11][19]  (.D(n5057), .SI(n8360), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[11][19] ), .QN(n8359));
   SDFFARX1 \key_mem_reg[12][19]  (.D(n5058), .SI(n8232), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[12][19] ), .QN(n8231));
   SDFFARX1 \key_mem_reg[13][19]  (.D(n5059), .SI(n8105), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7340), .Q(\key_mem[13][19] ), .QN(n8104));
   SDFFARX1 \key_mem_reg[14][19]  (.D(n5060), .SI(n7977), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[14][19] ), .QN(n7976));
   SDFFARX1 \prev_key1_reg_reg[18]  (.D(n5455), .SI(n7738), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(sboxw[18]), .QN(n7737));
   SDFFARX1 \prev_key0_reg_reg[18]  (.D(n5582), .SI(n7850), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(prev_key0_reg[18]), .QN(n7849));
   SDFFARX1 \key_mem_reg[0][18]  (.D(n5061), .SI(n9768), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[0][18] ), .QN(n9767));
   SDFFARX1 \key_mem_reg[1][18]  (.D(n5062), .SI(n9640), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[1][18] ), .QN(n9639));
   SDFFARX1 \key_mem_reg[2][18]  (.D(n5063), .SI(n9512), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[2][18] ), .QN(n9511));
   SDFFARX1 \key_mem_reg[3][18]  (.D(n5064), .SI(n9384), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[3][18] ), .QN(n9383));
   SDFFARX1 \key_mem_reg[4][18]  (.D(n5065), .SI(n9256), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[4][18] ), .QN(n9255));
   SDFFARX1 \key_mem_reg[5][18]  (.D(n5066), .SI(n9129), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[5][18] ), .QN(n9128));
   SDFFARX1 \key_mem_reg[6][18]  (.D(n5067), .SI(n9001), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[6][18] ), .QN(n9000));
   SDFFARX1 \key_mem_reg[7][18]  (.D(n5068), .SI(n8873), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[7][18] ), .QN(n8872));
   SDFFARX1 \key_mem_reg[8][18]  (.D(n5069), .SI(n8745), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7339), .Q(\key_mem[8][18] ), .QN(n8744));
   SDFFARX1 \key_mem_reg[9][18]  (.D(n5070), .SI(n8617), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[9][18] ), .QN(n8616));
   SDFFARX1 \key_mem_reg[10][18]  (.D(n5071), .SI(n8489), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[10][18] ), .QN(n8488));
   SDFFARX1 \key_mem_reg[11][18]  (.D(n5072), .SI(n8361), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[11][18] ), .QN(n8360));
   SDFFARX1 \key_mem_reg[12][18]  (.D(n5073), .SI(n8233), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[12][18] ), .QN(n8232));
   SDFFARX1 \key_mem_reg[13][18]  (.D(n5074), .SI(n8106), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[13][18] ), .QN(n8105));
   SDFFARX1 \key_mem_reg[14][18]  (.D(n5075), .SI(n7978), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[14][18] ), .QN(n7977));
   SDFFARX1 \prev_key1_reg_reg[17]  (.D(n5456), .SI(n7739), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(sboxw[17]), .QN(n7738));
   SDFFARX1 \prev_key0_reg_reg[17]  (.D(n5583), .SI(n7851), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(prev_key0_reg[17]), .QN(n7850));
   SDFFARX1 \key_mem_reg[0][17]  (.D(n5076), .SI(n9769), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[0][17] ), .QN(n9768));
   SDFFARX1 \key_mem_reg[1][17]  (.D(n5077), .SI(n9641), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[1][17] ), .QN(n9640));
   SDFFARX1 \key_mem_reg[2][17]  (.D(n5078), .SI(n9513), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[2][17] ), .QN(n9512));
   SDFFARX1 \key_mem_reg[3][17]  (.D(n5079), .SI(n9385), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7338), .Q(\key_mem[3][17] ), .QN(n9384));
   SDFFARX1 \key_mem_reg[4][17]  (.D(n5080), .SI(n9257), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[4][17] ), .QN(n9256));
   SDFFARX1 \key_mem_reg[5][17]  (.D(n5081), .SI(n9130), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[5][17] ), .QN(n9129));
   SDFFARX1 \key_mem_reg[6][17]  (.D(n5082), .SI(n9002), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[6][17] ), .QN(n9001));
   SDFFARX1 \key_mem_reg[7][17]  (.D(n5083), .SI(n8874), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[7][17] ), .QN(n8873));
   SDFFARX1 \key_mem_reg[8][17]  (.D(n5084), .SI(n8746), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[8][17] ), .QN(n8745));
   SDFFARX1 \key_mem_reg[9][17]  (.D(n5085), .SI(n8618), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[9][17] ), .QN(n8617));
   SDFFARX1 \key_mem_reg[10][17]  (.D(n5086), .SI(n8490), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[10][17] ), .QN(n8489));
   SDFFARX1 \key_mem_reg[11][17]  (.D(n5087), .SI(n8362), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[11][17] ), .QN(n8361));
   SDFFARX1 \key_mem_reg[12][17]  (.D(n5088), .SI(n8234), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[12][17] ), .QN(n8233));
   SDFFARX1 \key_mem_reg[13][17]  (.D(n5089), .SI(n8107), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[13][17] ), .QN(n8106));
   SDFFARX1 \key_mem_reg[14][17]  (.D(n5090), .SI(n7979), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(\key_mem[14][17] ), .QN(n7978));
   SDFFARX1 \prev_key1_reg_reg[16]  (.D(n5457), .SI(n7740), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7337), .Q(sboxw[16]), .QN(n7739));
   SDFFARX1 \prev_key0_reg_reg[16]  (.D(n5584), .SI(n7852), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(prev_key0_reg[16]), .QN(n7851));
   SDFFARX1 \key_mem_reg[0][16]  (.D(n5091), .SI(n9770), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[0][16] ), .QN(n9769));
   SDFFARX1 \key_mem_reg[1][16]  (.D(n5092), .SI(n9642), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[1][16] ), .QN(n9641));
   SDFFARX1 \key_mem_reg[2][16]  (.D(n5093), .SI(n9514), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[2][16] ), .QN(n9513));
   SDFFARX1 \key_mem_reg[3][16]  (.D(n5094), .SI(n9386), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[3][16] ), .QN(n9385));
   SDFFARX1 \key_mem_reg[4][16]  (.D(n5095), .SI(n9258), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[4][16] ), .QN(n9257));
   SDFFARX1 \key_mem_reg[5][16]  (.D(n5096), .SI(n9131), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[5][16] ), .QN(n9130));
   SDFFARX1 \key_mem_reg[6][16]  (.D(n5097), .SI(n9003), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[6][16] ), .QN(n9002));
   SDFFARX1 \key_mem_reg[7][16]  (.D(n5098), .SI(n8875), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[7][16] ), .QN(n8874));
   SDFFARX1 \key_mem_reg[8][16]  (.D(n5099), .SI(n8747), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[8][16] ), .QN(n8746));
   SDFFARX1 \key_mem_reg[9][16]  (.D(n5100), .SI(n8619), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[9][16] ), .QN(n8618));
   SDFFARX1 \key_mem_reg[10][16]  (.D(n5101), .SI(n8491), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7336), .Q(\key_mem[10][16] ), .QN(n8490));
   SDFFARX1 \key_mem_reg[11][16]  (.D(n5102), .SI(n8363), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[11][16] ), .QN(n8362));
   SDFFARX1 \key_mem_reg[12][16]  (.D(n5103), .SI(n8235), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[12][16] ), .QN(n8234));
   SDFFARX1 \key_mem_reg[13][16]  (.D(n5104), .SI(n8108), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[13][16] ), .QN(n8107));
   SDFFARX1 \key_mem_reg[14][16]  (.D(n5105), .SI(n7980), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[14][16] ), .QN(n7979));
   SDFFARX1 \prev_key1_reg_reg[15]  (.D(n5458), .SI(n7741), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(sboxw[15]), .QN(n7740));
   SDFFARX1 \prev_key0_reg_reg[15]  (.D(n5585), .SI(n7853), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(prev_key0_reg[15]), .QN(n7852));
   SDFFARX1 \key_mem_reg[0][15]  (.D(n5106), .SI(n9771), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[0][15] ), .QN(n9770));
   SDFFARX1 \key_mem_reg[1][15]  (.D(n5107), .SI(n9643), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[1][15] ), .QN(n9642));
   SDFFARX1 \key_mem_reg[2][15]  (.D(n5108), .SI(n9515), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[2][15] ), .QN(n9514));
   SDFFARX1 \key_mem_reg[3][15]  (.D(n5109), .SI(n9387), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[3][15] ), .QN(n9386));
   SDFFARX1 \key_mem_reg[4][15]  (.D(n5110), .SI(n9259), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[4][15] ), .QN(n9258));
   SDFFARX1 \key_mem_reg[5][15]  (.D(n5111), .SI(n9132), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7335), .Q(\key_mem[5][15] ), .QN(n9131));
   SDFFARX1 \key_mem_reg[6][15]  (.D(n5112), .SI(n9004), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[6][15] ), .QN(n9003));
   SDFFARX1 \key_mem_reg[7][15]  (.D(n5113), .SI(n8876), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[7][15] ), .QN(n8875));
   SDFFARX1 \key_mem_reg[8][15]  (.D(n5114), .SI(n8748), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[8][15] ), .QN(n8747));
   SDFFARX1 \key_mem_reg[9][15]  (.D(n5115), .SI(n8620), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[9][15] ), .QN(n8619));
   SDFFARX1 \key_mem_reg[10][15]  (.D(n5116), .SI(n8492), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[10][15] ), .QN(n8491));
   SDFFARX1 \key_mem_reg[11][15]  (.D(n5117), .SI(n8364), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[11][15] ), .QN(n8363));
   SDFFARX1 \key_mem_reg[12][15]  (.D(n5118), .SI(n8236), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[12][15] ), .QN(n8235));
   SDFFARX1 \key_mem_reg[13][15]  (.D(n5119), .SI(n8109), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[13][15] ), .QN(n8108));
   SDFFARX1 \key_mem_reg[14][15]  (.D(n5120), .SI(n7981), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[14][15] ), .QN(n7980));
   SDFFARX1 \prev_key1_reg_reg[14]  (.D(n5459), .SI(n7742), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(sboxw[14]), .QN(n7741));
   SDFFARX1 \prev_key0_reg_reg[14]  (.D(n5586), .SI(n7854), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(prev_key0_reg[14]), .QN(n7853));
   SDFFARX1 \key_mem_reg[0][14]  (.D(n5121), .SI(n9772), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7334), .Q(\key_mem[0][14] ), .QN(n9771));
   SDFFARX1 \key_mem_reg[1][14]  (.D(n5122), .SI(n9644), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[1][14] ), .QN(n9643));
   SDFFARX1 \key_mem_reg[2][14]  (.D(n5123), .SI(n9516), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[2][14] ), .QN(n9515));
   SDFFARX1 \key_mem_reg[3][14]  (.D(n5124), .SI(n9388), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[3][14] ), .QN(n9387));
   SDFFARX1 \key_mem_reg[4][14]  (.D(n5125), .SI(n9260), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[4][14] ), .QN(n9259));
   SDFFARX1 \key_mem_reg[5][14]  (.D(n5126), .SI(n9133), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[5][14] ), .QN(n9132));
   SDFFARX1 \key_mem_reg[6][14]  (.D(n5127), .SI(n9005), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[6][14] ), .QN(n9004));
   SDFFARX1 \key_mem_reg[7][14]  (.D(n5128), .SI(n8877), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[7][14] ), .QN(n8876));
   SDFFARX1 \key_mem_reg[8][14]  (.D(n5129), .SI(n8749), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[8][14] ), .QN(n8748));
   SDFFARX1 \key_mem_reg[9][14]  (.D(n5130), .SI(n8621), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[9][14] ), .QN(n8620));
   SDFFARX1 \key_mem_reg[10][14]  (.D(n5131), .SI(n8493), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[10][14] ), .QN(n8492));
   SDFFARX1 \key_mem_reg[11][14]  (.D(n5132), .SI(n8365), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[11][14] ), .QN(n8364));
   SDFFARX1 \key_mem_reg[12][14]  (.D(n5133), .SI(n8237), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7333), .Q(\key_mem[12][14] ), .QN(n8236));
   SDFFARX1 \key_mem_reg[13][14]  (.D(n5134), .SI(n8110), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[13][14] ), .QN(n8109));
   SDFFARX1 \key_mem_reg[14][14]  (.D(n5135), .SI(n7982), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[14][14] ), .QN(n7981));
   SDFFARX1 \prev_key1_reg_reg[13]  (.D(n5460), .SI(n7743), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(sboxw[13]), .QN(n7742));
   SDFFARX1 \prev_key0_reg_reg[13]  (.D(n5587), .SI(n7855), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(prev_key0_reg[13]), .QN(n7854));
   SDFFARX1 \key_mem_reg[0][13]  (.D(n5136), .SI(n9773), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[0][13] ), .QN(n9772));
   SDFFARX1 \key_mem_reg[1][13]  (.D(n5137), .SI(n9645), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[1][13] ), .QN(n9644));
   SDFFARX1 \key_mem_reg[2][13]  (.D(n5138), .SI(n9517), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[2][13] ), .QN(n9516));
   SDFFARX1 \key_mem_reg[3][13]  (.D(n5139), .SI(n9389), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[3][13] ), .QN(n9388));
   SDFFARX1 \key_mem_reg[4][13]  (.D(n5140), .SI(n9261), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[4][13] ), .QN(n9260));
   SDFFARX1 \key_mem_reg[5][13]  (.D(n5141), .SI(n9134), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[5][13] ), .QN(n9133));
   SDFFARX1 \key_mem_reg[6][13]  (.D(n5142), .SI(n9006), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[6][13] ), .QN(n9005));
   SDFFARX1 \key_mem_reg[7][13]  (.D(n5143), .SI(n8878), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7332), .Q(\key_mem[7][13] ), .QN(n8877));
   SDFFARX1 \key_mem_reg[8][13]  (.D(n5144), .SI(n8750), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[8][13] ), .QN(n8749));
   SDFFARX1 \key_mem_reg[9][13]  (.D(n5145), .SI(n8622), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[9][13] ), .QN(n8621));
   SDFFARX1 \key_mem_reg[10][13]  (.D(n5146), .SI(n8494), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[10][13] ), .QN(n8493));
   SDFFARX1 \key_mem_reg[11][13]  (.D(n5147), .SI(n8366), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[11][13] ), .QN(n8365));
   SDFFARX1 \key_mem_reg[12][13]  (.D(n5148), .SI(n8238), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[12][13] ), .QN(n8237));
   SDFFARX1 \key_mem_reg[13][13]  (.D(n5149), .SI(n8111), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[13][13] ), .QN(n8110));
   SDFFARX1 \key_mem_reg[14][13]  (.D(n5150), .SI(n7983), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[14][13] ), .QN(n7982));
   SDFFARX1 \prev_key1_reg_reg[12]  (.D(n5461), .SI(n7744), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(sboxw[12]), .QN(n7743));
   SDFFARX1 \prev_key0_reg_reg[12]  (.D(n5588), .SI(n7856), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(prev_key0_reg[12]), .QN(n7855));
   SDFFARX1 \key_mem_reg[0][12]  (.D(n5151), .SI(n9774), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[0][12] ), .QN(n9773));
   SDFFARX1 \key_mem_reg[1][12]  (.D(n5152), .SI(n9646), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[1][12] ), .QN(n9645));
   SDFFARX1 \key_mem_reg[2][12]  (.D(n5153), .SI(n9518), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7331), .Q(\key_mem[2][12] ), .QN(n9517));
   SDFFARX1 \key_mem_reg[3][12]  (.D(n5154), .SI(n9390), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[3][12] ), .QN(n9389));
   SDFFARX1 \key_mem_reg[4][12]  (.D(n5155), .SI(n9262), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[4][12] ), .QN(n9261));
   SDFFARX1 \key_mem_reg[5][12]  (.D(n5156), .SI(n9135), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[5][12] ), .QN(n9134));
   SDFFARX1 \key_mem_reg[6][12]  (.D(n5157), .SI(n9007), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[6][12] ), .QN(n9006));
   SDFFARX1 \key_mem_reg[7][12]  (.D(n5158), .SI(n8879), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[7][12] ), .QN(n8878));
   SDFFARX1 \key_mem_reg[8][12]  (.D(n5159), .SI(n8751), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[8][12] ), .QN(n8750));
   SDFFARX1 \key_mem_reg[9][12]  (.D(n5160), .SI(n8623), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[9][12] ), .QN(n8622));
   SDFFARX1 \key_mem_reg[10][12]  (.D(n5161), .SI(n8495), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[10][12] ), .QN(n8494));
   SDFFARX1 \key_mem_reg[11][12]  (.D(n5162), .SI(n8367), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[11][12] ), .QN(n8366));
   SDFFARX1 \key_mem_reg[12][12]  (.D(n5163), .SI(n8239), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[12][12] ), .QN(n8238));
   SDFFARX1 \key_mem_reg[13][12]  (.D(n5164), .SI(n8112), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[13][12] ), .QN(n8111));
   SDFFARX1 \key_mem_reg[14][12]  (.D(n5165), .SI(n7984), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7330), .Q(\key_mem[14][12] ), .QN(n7983));
   SDFFARX1 \prev_key1_reg_reg[11]  (.D(n5462), .SI(n7745), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(sboxw[11]), .QN(n7744));
   SDFFARX1 \prev_key0_reg_reg[11]  (.D(n5589), .SI(n7857), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(prev_key0_reg[11]), .QN(n7856));
   SDFFARX1 \key_mem_reg[0][11]  (.D(n5166), .SI(n9775), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[0][11] ), .QN(n9774));
   SDFFARX1 \key_mem_reg[1][11]  (.D(n5167), .SI(n9647), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[1][11] ), .QN(n9646));
   SDFFARX1 \key_mem_reg[2][11]  (.D(n5168), .SI(n9519), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[2][11] ), .QN(n9518));
   SDFFARX1 \key_mem_reg[3][11]  (.D(n5169), .SI(n9391), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[3][11] ), .QN(n9390));
   SDFFARX1 \key_mem_reg[4][11]  (.D(n5170), .SI(n9263), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[4][11] ), .QN(n9262));
   SDFFARX1 \key_mem_reg[5][11]  (.D(n5171), .SI(n9136), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[5][11] ), .QN(n9135));
   SDFFARX1 \key_mem_reg[6][11]  (.D(n5172), .SI(n9008), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[6][11] ), .QN(n9007));
   SDFFARX1 \key_mem_reg[7][11]  (.D(n5173), .SI(n8880), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[7][11] ), .QN(n8879));
   SDFFARX1 \key_mem_reg[8][11]  (.D(n5174), .SI(n8752), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[8][11] ), .QN(n8751));
   SDFFARX1 \key_mem_reg[9][11]  (.D(n5175), .SI(n8624), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7329), .Q(\key_mem[9][11] ), .QN(n8623));
   SDFFARX1 \key_mem_reg[10][11]  (.D(n5176), .SI(n8496), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[10][11] ), .QN(n8495));
   SDFFARX1 \key_mem_reg[11][11]  (.D(n5177), .SI(n8368), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[11][11] ), .QN(n8367));
   SDFFARX1 \key_mem_reg[12][11]  (.D(n5178), .SI(n8240), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[12][11] ), .QN(n8239));
   SDFFARX1 \key_mem_reg[13][11]  (.D(n5179), .SI(n8113), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[13][11] ), .QN(n8112));
   SDFFARX1 \key_mem_reg[14][11]  (.D(n5180), .SI(n7985), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[14][11] ), .QN(n7984));
   SDFFARX1 \prev_key1_reg_reg[10]  (.D(n5463), .SI(n7746), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(sboxw[10]), .QN(n7745));
   SDFFARX1 \prev_key0_reg_reg[10]  (.D(n5590), .SI(n7858), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(prev_key0_reg[10]), .QN(n7857));
   SDFFARX1 \key_mem_reg[0][10]  (.D(n5181), .SI(n9776), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[0][10] ), .QN(n9775));
   SDFFARX1 \key_mem_reg[1][10]  (.D(n5182), .SI(n9648), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[1][10] ), .QN(n9647));
   SDFFARX1 \key_mem_reg[2][10]  (.D(n5183), .SI(n9520), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[2][10] ), .QN(n9519));
   SDFFARX1 \key_mem_reg[3][10]  (.D(n5184), .SI(n9392), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[3][10] ), .QN(n9391));
   SDFFARX1 \key_mem_reg[4][10]  (.D(n5185), .SI(n9264), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7328), .Q(\key_mem[4][10] ), .QN(n9263));
   SDFFARX1 \key_mem_reg[5][10]  (.D(n5186), .SI(n9137), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[5][10] ), .QN(n9136));
   SDFFARX1 \key_mem_reg[6][10]  (.D(n5187), .SI(n9009), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[6][10] ), .QN(n9008));
   SDFFARX1 \key_mem_reg[7][10]  (.D(n5188), .SI(n8881), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[7][10] ), .QN(n8880));
   SDFFARX1 \key_mem_reg[8][10]  (.D(n5189), .SI(n8753), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[8][10] ), .QN(n8752));
   SDFFARX1 \key_mem_reg[9][10]  (.D(n5190), .SI(n8625), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[9][10] ), .QN(n8624));
   SDFFARX1 \key_mem_reg[10][10]  (.D(n5191), .SI(n8497), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[10][10] ), .QN(n8496));
   SDFFARX1 \key_mem_reg[11][10]  (.D(n5192), .SI(n8369), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[11][10] ), .QN(n8368));
   SDFFARX1 \key_mem_reg[12][10]  (.D(n5193), .SI(n8241), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[12][10] ), .QN(n8240));
   SDFFARX1 \key_mem_reg[13][10]  (.D(n5194), .SI(n8114), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[13][10] ), .QN(n8113));
   SDFFARX1 \key_mem_reg[14][10]  (.D(n5195), .SI(n7986), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(\key_mem[14][10] ), .QN(n7985));
   SDFFARX1 \prev_key1_reg_reg[9]  (.D(n5464), .SI(n7747), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(sboxw[9]), .QN(n7746));
   SDFFARX1 \prev_key0_reg_reg[9]  (.D(n5591), .SI(n7859), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7327), .Q(prev_key0_reg[9]), .QN(n7858));
   SDFFARX1 \key_mem_reg[0][9]  (.D(n5196), .SI(n9777), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[0][9] ), .QN(n9776));
   SDFFARX1 \key_mem_reg[1][9]  (.D(n5197), .SI(n9649), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[1][9] ), .QN(n9648));
   SDFFARX1 \key_mem_reg[2][9]  (.D(n5198), .SI(n9521), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[2][9] ), .QN(n9520));
   SDFFARX1 \key_mem_reg[3][9]  (.D(n5199), .SI(n9393), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[3][9] ), .QN(n9392));
   SDFFARX1 \key_mem_reg[4][9]  (.D(n5200), .SI(n9265), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[4][9] ), .QN(n9264));
   SDFFARX1 \key_mem_reg[5][9]  (.D(n5201), .SI(n9138), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[5][9] ), .QN(n9137));
   SDFFARX1 \key_mem_reg[6][9]  (.D(n5202), .SI(n9010), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[6][9] ), .QN(n9009));
   SDFFARX1 \key_mem_reg[7][9]  (.D(n5203), .SI(n8882), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[7][9] ), .QN(n8881));
   SDFFARX1 \key_mem_reg[8][9]  (.D(n5204), .SI(n8754), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[8][9] ), .QN(n8753));
   SDFFARX1 \key_mem_reg[9][9]  (.D(n5205), .SI(n8626), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[9][9] ), .QN(n8625));
   SDFFARX1 \key_mem_reg[10][9]  (.D(n5206), .SI(n8498), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[10][9] ), .QN(n8497));
   SDFFARX1 \key_mem_reg[11][9]  (.D(n5207), .SI(n8370), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7326), .Q(\key_mem[11][9] ), .QN(n8369));
   SDFFARX1 \key_mem_reg[12][9]  (.D(n5208), .SI(n8242), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[12][9] ), .QN(n8241));
   SDFFARX1 \key_mem_reg[13][9]  (.D(n5209), .SI(n8115), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[13][9] ), .QN(n8114));
   SDFFARX1 \key_mem_reg[14][9]  (.D(n5210), .SI(n7987), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[14][9] ), .QN(n7986));
   SDFFARX1 \prev_key1_reg_reg[8]  (.D(n5465), .SI(n7748), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(sboxw[8]), .QN(n7747));
   SDFFARX1 \prev_key0_reg_reg[8]  (.D(n5592), .SI(n7860), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(prev_key0_reg[8]), .QN(n7859));
   SDFFARX1 \key_mem_reg[0][8]  (.D(n5211), .SI(n9778), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[0][8] ), .QN(n9777));
   SDFFARX1 \key_mem_reg[1][8]  (.D(n5212), .SI(n9650), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[1][8] ), .QN(n9649));
   SDFFARX1 \key_mem_reg[2][8]  (.D(n5213), .SI(n9522), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[2][8] ), .QN(n9521));
   SDFFARX1 \key_mem_reg[3][8]  (.D(n5214), .SI(n9394), .SE(test_se_buf_net6), .CLK(
          clk_buf_net6), .RSTB(n7325), .Q(\key_mem[3][8] ), .QN(n9393));
   SDFFARX1 \key_mem_reg[4][8]  (.D(n5215), .SI(n9266), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7325), .Q(\key_mem[4][8] ), .QN(n9265));
   SDFFARX1 \key_mem_reg[5][8]  (.D(n5216), .SI(n9139), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7325), .Q(\key_mem[5][8] ), .QN(n9138));
   SDFFARX1 \key_mem_reg[6][8]  (.D(n5217), .SI(n9011), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7325), .Q(\key_mem[6][8] ), .QN(n9010));
   SDFFARX1 \key_mem_reg[7][8]  (.D(n5218), .SI(n8883), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[7][8] ), .QN(n8882));
   SDFFARX1 \key_mem_reg[8][8]  (.D(n5219), .SI(n8755), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[8][8] ), .QN(n8754));
   SDFFARX1 \key_mem_reg[9][8]  (.D(n5220), .SI(n8627), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[9][8] ), .QN(n8626));
   SDFFARX1 \key_mem_reg[10][8]  (.D(n5221), .SI(n8499), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[10][8] ), .QN(n8498));
   SDFFARX1 \key_mem_reg[11][8]  (.D(n5222), .SI(n8371), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[11][8] ), .QN(n8370));
   SDFFARX1 \key_mem_reg[12][8]  (.D(n5223), .SI(n8243), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[12][8] ), .QN(n8242));
   SDFFARX1 \key_mem_reg[13][8]  (.D(n5224), .SI(n8116), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[13][8] ), .QN(n8115));
   SDFFARX1 \key_mem_reg[14][8]  (.D(n5225), .SI(n7988), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[14][8] ), .QN(n7987));
   SDFFARX1 \prev_key1_reg_reg[7]  (.D(n5466), .SI(n7749), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(sboxw[7]), .QN(n7748));
   SDFFARX1 \prev_key0_reg_reg[7]  (.D(n5593), .SI(n7861), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(prev_key0_reg[7]), .QN(n7860));
   SDFFARX1 \key_mem_reg[0][7]  (.D(n5226), .SI(n9779), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[0][7] ), .QN(n9778));
   SDFFARX1 \key_mem_reg[1][7]  (.D(n5227), .SI(n9651), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7324), .Q(\key_mem[1][7] ), .QN(n9650));
   SDFFARX1 \key_mem_reg[2][7]  (.D(n5228), .SI(n9523), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[2][7] ), .QN(n9522));
   SDFFARX1 \key_mem_reg[3][7]  (.D(n5229), .SI(n9395), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[3][7] ), .QN(n9394));
   SDFFARX1 \key_mem_reg[4][7]  (.D(n5230), .SI(n9267), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[4][7] ), .QN(n9266));
   SDFFARX1 \key_mem_reg[5][7]  (.D(n5231), .SI(n9140), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[5][7] ), .QN(n9139));
   SDFFARX1 \key_mem_reg[6][7]  (.D(n5232), .SI(n9012), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[6][7] ), .QN(n9011));
   SDFFARX1 \key_mem_reg[7][7]  (.D(n5233), .SI(n8884), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[7][7] ), .QN(n8883));
   SDFFARX1 \key_mem_reg[8][7]  (.D(n5234), .SI(n8756), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[8][7] ), .QN(n8755));
   SDFFARX1 \key_mem_reg[9][7]  (.D(n5235), .SI(n8628), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[9][7] ), .QN(n8627));
   SDFFARX1 \key_mem_reg[10][7]  (.D(n5236), .SI(n8500), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[10][7] ), .QN(n8499));
   SDFFARX1 \key_mem_reg[11][7]  (.D(n5237), .SI(n8372), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[11][7] ), .QN(n8371));
   SDFFARX1 \key_mem_reg[12][7]  (.D(n5238), .SI(n8244), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[12][7] ), .QN(n8243));
   SDFFARX1 \key_mem_reg[13][7]  (.D(n5239), .SI(n8117), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7323), .Q(\key_mem[13][7] ), .QN(n8116));
   SDFFARX1 \key_mem_reg[14][7]  (.D(n5240), .SI(n7989), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[14][7] ), .QN(n7988));
   SDFFARX1 \prev_key1_reg_reg[6]  (.D(n5467), .SI(n7750), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(sboxw[6]), .QN(n7749));
   SDFFARX1 \prev_key0_reg_reg[6]  (.D(n5594), .SI(n7862), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(prev_key0_reg[6]), .QN(n7861));
   SDFFARX1 \key_mem_reg[0][6]  (.D(n5241), .SI(n9780), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[0][6] ), .QN(n9779));
   SDFFARX1 \key_mem_reg[1][6]  (.D(n5242), .SI(n9652), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[1][6] ), .QN(n9651));
   SDFFARX1 \key_mem_reg[2][6]  (.D(n5243), .SI(n9524), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[2][6] ), .QN(n9523));
   SDFFARX1 \key_mem_reg[3][6]  (.D(n5244), .SI(n9396), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[3][6] ), .QN(n9395));
   SDFFARX1 \key_mem_reg[4][6]  (.D(n5245), .SI(n9268), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[4][6] ), .QN(n9267));
   SDFFARX1 \key_mem_reg[5][6]  (.D(n5246), .SI(n9141), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[5][6] ), .QN(n9140));
   SDFFARX1 \key_mem_reg[6][6]  (.D(n5247), .SI(n9013), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[6][6] ), .QN(n9012));
   SDFFARX1 \key_mem_reg[7][6]  (.D(n5248), .SI(n8885), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[7][6] ), .QN(n8884));
   SDFFARX1 \key_mem_reg[8][6]  (.D(n5249), .SI(n8757), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7322), .Q(\key_mem[8][6] ), .QN(n8756));
   SDFFARX1 \key_mem_reg[9][6]  (.D(n5250), .SI(n8629), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[9][6] ), .QN(n8628));
   SDFFARX1 \key_mem_reg[10][6]  (.D(n5251), .SI(n8501), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[10][6] ), .QN(n8500));
   SDFFARX1 \key_mem_reg[11][6]  (.D(n5252), .SI(n8373), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[11][6] ), .QN(n8372));
   SDFFARX1 \key_mem_reg[12][6]  (.D(n5253), .SI(n8245), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[12][6] ), .QN(n8244));
   SDFFARX1 \key_mem_reg[13][6]  (.D(n5254), .SI(n8118), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[13][6] ), .QN(n8117));
   SDFFARX1 \key_mem_reg[14][6]  (.D(n5255), .SI(n7990), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[14][6] ), .QN(n7989));
   SDFFARX1 \prev_key1_reg_reg[5]  (.D(n5468), .SI(n7751), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(sboxw[5]), .QN(n7750));
   SDFFARX1 \prev_key0_reg_reg[5]  (.D(n5595), .SI(n7863), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(prev_key0_reg[5]), .QN(n7862));
   SDFFARX1 \key_mem_reg[0][5]  (.D(n5256), .SI(n9781), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[0][5] ), .QN(n9780));
   SDFFARX1 \key_mem_reg[1][5]  (.D(n5257), .SI(n9653), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[1][5] ), .QN(n9652));
   SDFFARX1 \key_mem_reg[2][5]  (.D(n5258), .SI(n9525), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[2][5] ), .QN(n9524));
   SDFFARX1 \key_mem_reg[3][5]  (.D(n5259), .SI(n9397), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7321), .Q(\key_mem[3][5] ), .QN(n9396));
   SDFFARX1 \key_mem_reg[4][5]  (.D(n5260), .SI(n9269), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[4][5] ), .QN(n9268));
   SDFFARX1 \key_mem_reg[5][5]  (.D(n5261), .SI(n9142), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[5][5] ), .QN(n9141));
   SDFFARX1 \key_mem_reg[6][5]  (.D(n5262), .SI(n9014), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[6][5] ), .QN(n9013));
   SDFFARX1 \key_mem_reg[7][5]  (.D(n5263), .SI(n8886), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[7][5] ), .QN(n8885));
   SDFFARX1 \key_mem_reg[8][5]  (.D(n5264), .SI(n8758), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[8][5] ), .QN(n8757));
   SDFFARX1 \key_mem_reg[9][5]  (.D(n5265), .SI(n8630), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[9][5] ), .QN(n8629));
   SDFFARX1 \key_mem_reg[10][5]  (.D(n5266), .SI(n8502), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[10][5] ), .QN(n8501));
   SDFFARX1 \key_mem_reg[11][5]  (.D(n5267), .SI(n8374), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[11][5] ), .QN(n8373));
   SDFFARX1 \key_mem_reg[12][5]  (.D(n5268), .SI(n8246), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[12][5] ), .QN(n8245));
   SDFFARX1 \key_mem_reg[13][5]  (.D(n5269), .SI(n8119), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[13][5] ), .QN(n8118));
   SDFFARX1 \key_mem_reg[14][5]  (.D(n5270), .SI(n7991), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(\key_mem[14][5] ), .QN(n7990));
   SDFFARX1 \prev_key1_reg_reg[4]  (.D(n5469), .SI(n7752), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7320), .Q(sboxw[4]), .QN(n7751));
   SDFFARX1 \prev_key0_reg_reg[4]  (.D(n5596), .SI(n7864), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(prev_key0_reg[4]), .QN(n7863));
   SDFFARX1 \key_mem_reg[0][4]  (.D(n5271), .SI(n9782), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[0][4] ), .QN(n9781));
   SDFFARX1 \key_mem_reg[1][4]  (.D(n5272), .SI(n9654), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[1][4] ), .QN(n9653));
   SDFFARX1 \key_mem_reg[2][4]  (.D(n5273), .SI(n9526), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[2][4] ), .QN(n9525));
   SDFFARX1 \key_mem_reg[3][4]  (.D(n5274), .SI(n9398), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[3][4] ), .QN(n9397));
   SDFFARX1 \key_mem_reg[4][4]  (.D(n5275), .SI(n9270), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[4][4] ), .QN(n9269));
   SDFFARX1 \key_mem_reg[5][4]  (.D(n5276), .SI(n9143), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[5][4] ), .QN(n9142));
   SDFFARX1 \key_mem_reg[6][4]  (.D(n5277), .SI(n9015), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[6][4] ), .QN(n9014));
   SDFFARX1 \key_mem_reg[7][4]  (.D(n5278), .SI(n8887), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[7][4] ), .QN(n8886));
   SDFFARX1 \key_mem_reg[8][4]  (.D(n5279), .SI(n8759), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[8][4] ), .QN(n8758));
   SDFFARX1 \key_mem_reg[9][4]  (.D(n5280), .SI(n8631), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[9][4] ), .QN(n8630));
   SDFFARX1 \key_mem_reg[10][4]  (.D(n5281), .SI(n8503), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7319), .Q(\key_mem[10][4] ), .QN(n8502));
   SDFFARX1 \key_mem_reg[11][4]  (.D(n5282), .SI(n8375), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[11][4] ), .QN(n8374));
   SDFFARX1 \key_mem_reg[12][4]  (.D(n5283), .SI(n8247), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[12][4] ), .QN(n8246));
   SDFFARX1 \key_mem_reg[13][4]  (.D(n5284), .SI(n8120), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[13][4] ), .QN(n8119));
   SDFFARX1 \key_mem_reg[14][4]  (.D(n5285), .SI(n7992), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[14][4] ), .QN(n7991));
   SDFFARX1 \prev_key1_reg_reg[3]  (.D(n5470), .SI(n7753), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(sboxw[3]), .QN(n7752));
   SDFFARX1 \prev_key0_reg_reg[3]  (.D(n5597), .SI(n7865), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(prev_key0_reg[3]), .QN(n7864));
   SDFFARX1 \key_mem_reg[0][3]  (.D(n5286), .SI(n9783), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[0][3] ), .QN(n9782));
   SDFFARX1 \key_mem_reg[1][3]  (.D(n5287), .SI(n9655), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[1][3] ), .QN(n9654));
   SDFFARX1 \key_mem_reg[2][3]  (.D(n5288), .SI(n9527), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[2][3] ), .QN(n9526));
   SDFFARX1 \key_mem_reg[3][3]  (.D(n5289), .SI(n9399), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[3][3] ), .QN(n9398));
   SDFFARX1 \key_mem_reg[4][3]  (.D(n5290), .SI(n9271), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[4][3] ), .QN(n9270));
   SDFFARX1 \key_mem_reg[5][3]  (.D(n5291), .SI(n9144), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7318), .Q(\key_mem[5][3] ), .QN(n9143));
   SDFFARX1 \key_mem_reg[6][3]  (.D(n5292), .SI(n9016), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[6][3] ), .QN(n9015));
   SDFFARX1 \key_mem_reg[7][3]  (.D(n5293), .SI(n8888), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[7][3] ), .QN(n8887));
   SDFFARX1 \key_mem_reg[8][3]  (.D(n5294), .SI(n8760), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[8][3] ), .QN(n8759));
   SDFFARX1 \key_mem_reg[9][3]  (.D(n5295), .SI(n8632), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[9][3] ), .QN(n8631));
   SDFFARX1 \key_mem_reg[10][3]  (.D(n5296), .SI(n8504), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[10][3] ), .QN(n8503));
   SDFFARX1 \key_mem_reg[11][3]  (.D(n5297), .SI(n8376), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[11][3] ), .QN(n8375));
   SDFFARX1 \key_mem_reg[12][3]  (.D(n5298), .SI(n8248), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[12][3] ), .QN(n8247));
   SDFFARX1 \key_mem_reg[13][3]  (.D(n5299), .SI(n8121), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[13][3] ), .QN(n8120));
   SDFFARX1 \key_mem_reg[14][3]  (.D(n5300), .SI(n7993), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[14][3] ), .QN(n7992));
   SDFFARX1 \prev_key1_reg_reg[2]  (.D(n5471), .SI(n7754), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(sboxw[2]), .QN(n7753));
   SDFFARX1 \prev_key0_reg_reg[2]  (.D(n5598), .SI(n7866), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(prev_key0_reg[2]), .QN(n7865));
   SDFFARX1 \key_mem_reg[0][2]  (.D(n5301), .SI(n9784), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7317), .Q(\key_mem[0][2] ), .QN(n9783));
   SDFFARX1 \key_mem_reg[1][2]  (.D(n5302), .SI(n9656), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[1][2] ), .QN(n9655));
   SDFFARX1 \key_mem_reg[2][2]  (.D(n5303), .SI(n9528), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[2][2] ), .QN(n9527));
   SDFFARX1 \key_mem_reg[3][2]  (.D(n5304), .SI(n9400), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[3][2] ), .QN(n9399));
   SDFFARX1 \key_mem_reg[4][2]  (.D(n5305), .SI(n9272), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[4][2] ), .QN(n9271));
   SDFFARX1 \key_mem_reg[5][2]  (.D(n5306), .SI(n9145), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[5][2] ), .QN(n9144));
   SDFFARX1 \key_mem_reg[6][2]  (.D(n5307), .SI(n9017), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[6][2] ), .QN(n9016));
   SDFFARX1 \key_mem_reg[7][2]  (.D(n5308), .SI(n8889), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[7][2] ), .QN(n8888));
   SDFFARX1 \key_mem_reg[8][2]  (.D(n5309), .SI(n8761), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[8][2] ), .QN(n8760));
   SDFFARX1 \key_mem_reg[9][2]  (.D(n5310), .SI(n8633), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[9][2] ), .QN(n8632));
   SDFFARX1 \key_mem_reg[10][2]  (.D(n5311), .SI(n8505), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[10][2] ), .QN(n8504));
   SDFFARX1 \key_mem_reg[11][2]  (.D(n5312), .SI(n8377), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[11][2] ), .QN(n8376));
   SDFFARX1 \key_mem_reg[12][2]  (.D(n5313), .SI(n8249), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7316), .Q(\key_mem[12][2] ), .QN(n8248));
   SDFFARX1 \key_mem_reg[13][2]  (.D(n5314), .SI(n8122), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[13][2] ), .QN(n8121));
   SDFFARX1 \key_mem_reg[14][2]  (.D(n5315), .SI(n7994), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[14][2] ), .QN(n7993));
   SDFFARX1 \prev_key1_reg_reg[1]  (.D(n5472), .SI(n7755), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(sboxw[1]), .QN(n7754));
   SDFFARX1 \prev_key0_reg_reg[1]  (.D(n5599), .SI(n7867), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(prev_key0_reg[1]), .QN(n7866));
   SDFFARX1 \key_mem_reg[0][1]  (.D(n5316), .SI(n9785), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[0][1] ), .QN(n9784));
   SDFFARX1 \key_mem_reg[1][1]  (.D(n5317), .SI(n9657), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[1][1] ), .QN(n9656));
   SDFFARX1 \key_mem_reg[2][1]  (.D(n5318), .SI(n9529), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[2][1] ), .QN(n9528));
   SDFFARX1 \key_mem_reg[3][1]  (.D(n5319), .SI(n9401), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[3][1] ), .QN(n9400));
   SDFFARX1 \key_mem_reg[4][1]  (.D(n5320), .SI(n9273), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[4][1] ), .QN(n9272));
   SDFFARX1 \key_mem_reg[5][1]  (.D(n5321), .SI(n9146), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[5][1] ), .QN(n9145));
   SDFFARX1 \key_mem_reg[6][1]  (.D(n5322), .SI(n9018), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[6][1] ), .QN(n9017));
   SDFFARX1 \key_mem_reg[7][1]  (.D(n5323), .SI(n8890), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7315), .Q(\key_mem[7][1] ), .QN(n8889));
   SDFFARX1 \key_mem_reg[8][1]  (.D(n5324), .SI(n8762), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[8][1] ), .QN(n8761));
   SDFFARX1 \key_mem_reg[9][1]  (.D(n5325), .SI(n8634), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[9][1] ), .QN(n8633));
   SDFFARX1 \key_mem_reg[10][1]  (.D(n5326), .SI(n8506), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[10][1] ), .QN(n8505));
   SDFFARX1 \key_mem_reg[11][1]  (.D(n5327), .SI(n8378), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[11][1] ), .QN(n8377));
   SDFFARX1 \key_mem_reg[12][1]  (.D(n5328), .SI(n8250), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[12][1] ), .QN(n8249));
   SDFFARX1 \key_mem_reg[13][1]  (.D(n5329), .SI(n8123), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[13][1] ), .QN(n8122));
   SDFFARX1 \key_mem_reg[14][1]  (.D(n5330), .SI(n7995), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[14][1] ), .QN(n7994));
   SDFFARX1 \prev_key1_reg_reg[0]  (.D(n5601), .SI(prev_key0_reg[127]), .SE(
          test_se_buf_net7), .CLK(clk_buf_net7), .RSTB(n7314), .Q(sboxw[0]), .QN(n7755));
   SDFFARX1 \prev_key0_reg_reg[0]  (.D(n5600), .SI(n7868), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(prev_key0_reg[0]), .QN(n7867));
   SDFFARX1 \key_mem_reg[0][0]  (.D(n5331), .SI(n2242), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[0][0] ), .QN(n9785));
   SDFFARX1 \key_mem_reg[1][0]  (.D(n5332), .SI(n9658), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[1][0] ), .QN(n9657));
   SDFFARX1 \key_mem_reg[2][0]  (.D(n5333), .SI(n9530), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7314), .Q(\key_mem[2][0] ), .QN(n9529));
   SDFFARX1 \key_mem_reg[3][0]  (.D(n5334), .SI(n9402), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[3][0] ), .QN(n9401));
   SDFFARX1 \key_mem_reg[4][0]  (.D(n5335), .SI(n9274), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[4][0] ), .QN(n9273));
   SDFFARX1 \key_mem_reg[5][0]  (.D(n5336), .SI(n9147), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[5][0] ), .QN(n9146));
   SDFFARX1 \key_mem_reg[6][0]  (.D(n5337), .SI(n9019), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[6][0] ), .QN(n9018));
   SDFFARX1 \key_mem_reg[7][0]  (.D(n5338), .SI(n8891), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[7][0] ), .QN(n8890));
   SDFFARX1 \key_mem_reg[8][0]  (.D(n5339), .SI(n8763), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[8][0] ), .QN(n8762));
   SDFFARX1 \key_mem_reg[9][0]  (.D(n5340), .SI(n8635), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[9][0] ), .QN(n8634));
   SDFFARX1 \key_mem_reg[10][0]  (.D(n5341), .SI(n8507), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[10][0] ), .QN(n8506));
   SDFFARX1 \key_mem_reg[11][0]  (.D(n5342), .SI(n8379), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[11][0] ), .QN(n8378));
   SDFFARX1 \key_mem_reg[12][0]  (.D(n5343), .SI(n8251), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[12][0] ), .QN(n8250));
   SDFFARX1 \key_mem_reg[13][0]  (.D(n5344), .SI(n8124), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[13][0] ), .QN(n8123));
   SDFFARX1 \key_mem_reg[14][0]  (.D(n5345), .SI(n7996), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7313), .Q(\key_mem[14][0] ), .QN(n7995));
   AO22X1 U2406 (.IN1(n7299), .IN2(n2277), .IN3(\key_mem[0][127] ), .IN4(n6938), .Q(n3426)
          );
   AO22X1 U2407 (.IN1(n6809), .IN2(n2277), .IN3(\key_mem[1][127] ), .IN4(n6825), .Q(n3427)
          );
   AO22X1 U2408 (.IN1(n6853), .IN2(n2277), .IN3(\key_mem[2][127] ), .IN4(n6848), .Q(n3428)
          );
   AO22X1 U2409 (.IN1(n6869), .IN2(n2277), .IN3(\key_mem[3][127] ), .IN4(n6864), .Q(n3429)
          );
   AO22X1 U2410 (.IN1(n6887), .IN2(n2277), .IN3(\key_mem[4][127] ), .IN4(n6923), .Q(n3430)
          );
   AO22X1 U2411 (.IN1(n6973), .IN2(n2277), .IN3(\key_mem[5][127] ), .IN4(n7018), .Q(n3431)
          );
   AO22X1 U2412 (.IN1(n7262), .IN2(n2277), .IN3(\key_mem[6][127] ), .IN4(n7257), .Q(n3432)
          );
   AO22X1 U2413 (.IN1(n7014), .IN2(n2277), .IN3(\key_mem[7][127] ), .IN4(n7237), .Q(n3433)
          );
   AO22X1 U2414 (.IN1(n6750), .IN2(n2277), .IN3(\key_mem[8][127] ), .IN4(n6747), .Q(n3434)
          );
   AO22X1 U2415 (.IN1(n6975), .IN2(n2277), .IN3(\key_mem[9][127] ), .IN4(n7217), .Q(n3435)
          );
   AO22X1 U2416 (.IN1(n6797), .IN2(n2277), .IN3(\key_mem[10][127] ), .IN4(n6794), .Q(n3436)
          );
   AO22X1 U2417 (.IN1(n6977), .IN2(n2277), .IN3(\key_mem[11][127] ), .IN4(n7193), .Q(n3437)
          );
   AO22X1 U2418 (.IN1(n6840), .IN2(n2277), .IN3(\key_mem[12][127] ), .IN4(n7000), .Q(n3438)
          );
   AO22X1 U2419 (.IN1(n6979), .IN2(n2277), .IN3(\key_mem[13][127] ), .IN4(n7172), .Q(n3439)
          );
   AO22X1 U2420 (.IN1(n7162), .IN2(n2277), .IN3(\key_mem[14][127] ), .IN4(n7156), .Q(n3440)
          );
   AO222X1 U2422 (.IN1(n7118), .IN2(n2296), .IN3(key[127]), .IN4(n7071), .IN5(n7038), .IN6(
          n2299), .Q(n2294));
   AO22X1 U2423 (.IN1(n7299), .IN2(n2300), .IN3(\key_mem[0][126] ), .IN4(n6938), .Q(n3441)
          );
   AO22X1 U2424 (.IN1(n6811), .IN2(n2300), .IN3(\key_mem[1][126] ), .IN4(n6821), .Q(n3442)
          );
   AO22X1 U2425 (.IN1(n6856), .IN2(n2300), .IN3(\key_mem[2][126] ), .IN4(n6849), .Q(n3443)
          );
   AO22X1 U2426 (.IN1(n6989), .IN2(n2300), .IN3(\key_mem[3][126] ), .IN4(n6877), .Q(n3444)
          );
   AO22X1 U2427 (.IN1(n6888), .IN2(n2300), .IN3(\key_mem[4][126] ), .IN4(n6923), .Q(n3445)
          );
   AO22X1 U2428 (.IN1(n7274), .IN2(n2300), .IN3(\key_mem[5][126] ), .IN4(n7270), .Q(n3446)
          );
   AO22X1 U2429 (.IN1(n7016), .IN2(n2300), .IN3(\key_mem[6][126] ), .IN4(n7254), .Q(n3447)
          );
   AO22X1 U2430 (.IN1(n7246), .IN2(n2300), .IN3(\key_mem[7][126] ), .IN4(n2284), .Q(n3448)
          );
   AO22X1 U2431 (.IN1(n6751), .IN2(n2300), .IN3(\key_mem[8][126] ), .IN4(n6715), .Q(n3449)
          );
   AO22X1 U2432 (.IN1(n7218), .IN2(n2300), .IN3(\key_mem[9][126] ), .IN4(n7226), .Q(n3450)
          );
   AO22X1 U2433 (.IN1(n6798), .IN2(n2300), .IN3(\key_mem[10][126] ), .IN4(n6762), .Q(n3451)
          );
   AO22X1 U2434 (.IN1(n7194), .IN2(n2300), .IN3(\key_mem[11][126] ), .IN4(n7202), .Q(n3452)
          );
   AO22X1 U2435 (.IN1(n7186), .IN2(n2300), .IN3(\key_mem[12][126] ), .IN4(n6828), .Q(n3453)
          );
   AO22X1 U2436 (.IN1(n7173), .IN2(n2300), .IN3(\key_mem[13][126] ), .IN4(n7181), .Q(n3454)
          );
   AO22X1 U2437 (.IN1(n7161), .IN2(n2300), .IN3(\key_mem[14][126] ), .IN4(n7157), .Q(n3455)
          );
   AO221X1 U2438 (.IN1(n7126), .IN2(n2301), .IN3(key[254]), .IN4(n7312), .IN5(n2302), .Q(
          n2300));
   AO222X1 U2439 (.IN1(n7118), .IN2(n2303), .IN3(key[126]), .IN4(n7071), .IN5(n7038), .IN6(
          n2304), .Q(n2302));
   AO22X1 U2440 (.IN1(n7292), .IN2(n2305), .IN3(\key_mem[0][125] ), .IN4(n6938), .Q(n3456)
          );
   AO22X1 U2441 (.IN1(n6812), .IN2(n2305), .IN3(\key_mem[1][125] ), .IN4(n6815), .Q(n3457)
          );
   AO22X1 U2442 (.IN1(n6858), .IN2(n2305), .IN3(\key_mem[2][125] ), .IN4(n6844), .Q(n3458)
          );
   AO22X1 U2443 (.IN1(n6870), .IN2(n2305), .IN3(\key_mem[3][125] ), .IN4(n6860), .Q(n3459)
          );
   AO22X1 U2444 (.IN1(n6922), .IN2(n2305), .IN3(\key_mem[4][125] ), .IN4(n7284), .Q(n3460)
          );
   AO22X1 U2445 (.IN1(n7279), .IN2(n2305), .IN3(\key_mem[5][125] ), .IN4(n7268), .Q(n3461)
          );
   AO22X1 U2446 (.IN1(n7263), .IN2(n2305), .IN3(\key_mem[6][125] ), .IN4(n7255), .Q(n3462)
          );
   AO22X1 U2447 (.IN1(n7246), .IN2(n2305), .IN3(\key_mem[7][125] ), .IN4(n7012), .Q(n3463)
          );
   AO22X1 U2448 (.IN1(n6752), .IN2(n2305), .IN3(\key_mem[8][125] ), .IN4(n7228), .Q(n3464)
          );
   AO22X1 U2449 (.IN1(n7223), .IN2(n2305), .IN3(\key_mem[9][125] ), .IN4(n7217), .Q(n3465)
          );
   AO22X1 U2450 (.IN1(n6799), .IN2(n2305), .IN3(\key_mem[10][125] ), .IN4(n7204), .Q(n3466)
          );
   AO22X1 U2451 (.IN1(n7199), .IN2(n2305), .IN3(\key_mem[11][125] ), .IN4(n7193), .Q(n3467)
          );
   AO22X1 U2452 (.IN1(n6832), .IN2(n2305), .IN3(\key_mem[12][125] ), .IN4(n7185), .Q(n3468)
          );
   AO22X1 U2453 (.IN1(n7178), .IN2(n2305), .IN3(\key_mem[13][125] ), .IN4(n7172), .Q(n3469)
          );
   AO22X1 U2454 (.IN1(n7158), .IN2(n2305), .IN3(\key_mem[14][125] ), .IN4(n7154), .Q(n3470)
          );
   AO222X1 U2456 (.IN1(n7118), .IN2(n2308), .IN3(key[125]), .IN4(n7071), .IN5(n7038), .IN6(
          n2309), .Q(n2307));
   AO22X1 U2457 (.IN1(n7297), .IN2(n2310), .IN3(\key_mem[0][124] ), .IN4(n6938), .Q(n3471)
          );
   AO22X1 U2458 (.IN1(n6813), .IN2(n2310), .IN3(\key_mem[1][124] ), .IN4(n6817), .Q(n3472)
          );
   AO22X1 U2459 (.IN1(n6857), .IN2(n2310), .IN3(\key_mem[2][124] ), .IN4(n6850), .Q(n3473)
          );
   AO22X1 U2460 (.IN1(n6874), .IN2(n2310), .IN3(\key_mem[3][124] ), .IN4(n6868), .Q(n3474)
          );
   AO22X1 U2461 (.IN1(n6922), .IN2(n2310), .IN3(\key_mem[4][124] ), .IN4(n7021), .Q(n3475)
          );
   AO22X1 U2462 (.IN1(n7276), .IN2(n2310), .IN3(\key_mem[5][124] ), .IN4(n7269), .Q(n3476)
          );
   AO22X1 U2463 (.IN1(n7263), .IN2(n2310), .IN3(\key_mem[6][124] ), .IN4(n7252), .Q(n3477)
          );
   AO22X1 U2464 (.IN1(n7245), .IN2(n2310), .IN3(\key_mem[7][124] ), .IN4(n7243), .Q(n3478)
          );
   AO22X1 U2465 (.IN1(n6754), .IN2(n2310), .IN3(\key_mem[8][124] ), .IN4(n6721), .Q(n3479)
          );
   AO22X1 U2466 (.IN1(n7220), .IN2(n2310), .IN3(\key_mem[9][124] ), .IN4(n7215), .Q(n3480)
          );
   AO22X1 U2467 (.IN1(n6801), .IN2(n2310), .IN3(\key_mem[10][124] ), .IN4(n6768), .Q(n3481)
          );
   AO22X1 U2468 (.IN1(n7196), .IN2(n2310), .IN3(\key_mem[11][124] ), .IN4(n7191), .Q(n3482)
          );
   AO22X1 U2469 (.IN1(n6835), .IN2(n2310), .IN3(\key_mem[12][124] ), .IN4(n6836), .Q(n3483)
          );
   AO22X1 U2470 (.IN1(n7175), .IN2(n2310), .IN3(\key_mem[13][124] ), .IN4(n7170), .Q(n3484)
          );
   AO22X1 U2471 (.IN1(n6995), .IN2(n2310), .IN3(\key_mem[14][124] ), .IN4(n7155), .Q(n3485)
          );
   AO222X1 U2473 (.IN1(n7118), .IN2(n2313), .IN3(key[124]), .IN4(n7071), .IN5(n7038), .IN6(
          n2314), .Q(n2312));
   AO22X1 U2474 (.IN1(n7292), .IN2(n2315), .IN3(\key_mem[0][123] ), .IN4(n6938), .Q(n3486)
          );
   AO22X1 U2475 (.IN1(n6809), .IN2(n2315), .IN3(\key_mem[1][123] ), .IN4(n6819), .Q(n3487)
          );
   AO22X1 U2476 (.IN1(n6988), .IN2(n2315), .IN3(\key_mem[2][123] ), .IN4(n6847), .Q(n3488)
          );
   AO22X1 U2477 (.IN1(n6875), .IN2(n2315), .IN3(\key_mem[3][123] ), .IN4(n6868), .Q(n3489)
          );
   AO22X1 U2478 (.IN1(n7286), .IN2(n2315), .IN3(\key_mem[4][123] ), .IN4(n7284), .Q(n3490)
          );
   AO22X1 U2479 (.IN1(n7277), .IN2(n2315), .IN3(\key_mem[5][123] ), .IN4(n7268), .Q(n3491)
          );
   AO22X1 U2480 (.IN1(n7263), .IN2(n2315), .IN3(\key_mem[6][123] ), .IN4(n7253), .Q(n3492)
          );
   AO22X1 U2481 (.IN1(n7244), .IN2(n2315), .IN3(\key_mem[7][123] ), .IN4(n7235), .Q(n3493)
          );
   AO22X1 U2482 (.IN1(n6751), .IN2(n2315), .IN3(\key_mem[8][123] ), .IN4(n6724), .Q(n3494)
          );
   AO22X1 U2483 (.IN1(n7221), .IN2(n2315), .IN3(\key_mem[9][123] ), .IN4(n7216), .Q(n3495)
          );
   AO22X1 U2484 (.IN1(n6798), .IN2(n2315), .IN3(\key_mem[10][123] ), .IN4(n6771), .Q(n3496)
          );
   AO22X1 U2485 (.IN1(n7197), .IN2(n2315), .IN3(\key_mem[11][123] ), .IN4(n7192), .Q(n3497)
          );
   AO22X1 U2486 (.IN1(n7001), .IN2(n2315), .IN3(\key_mem[12][123] ), .IN4(n6841), .Q(n3498)
          );
   AO22X1 U2487 (.IN1(n7176), .IN2(n2315), .IN3(\key_mem[13][123] ), .IN4(n7171), .Q(n3499)
          );
   AO22X1 U2488 (.IN1(n7162), .IN2(n2315), .IN3(\key_mem[14][123] ), .IN4(n7147), .Q(n3500)
          );
   AO221X1 U2489 (.IN1(n7126), .IN2(n2316), .IN3(key[251]), .IN4(n7306), .IN5(n2317), .Q(
          n2315));
   AO222X1 U2490 (.IN1(n7118), .IN2(n2318), .IN3(key[123]), .IN4(n7071), .IN5(n7038), .IN6(
          n2319), .Q(n2317));
   AO22X1 U2491 (.IN1(n7301), .IN2(n2320), .IN3(\key_mem[0][122] ), .IN4(n6938), .Q(n3501)
          );
   AO22X1 U2492 (.IN1(n6926), .IN2(n2320), .IN3(\key_mem[1][122] ), .IN4(n6820), .Q(n3502)
          );
   AO22X1 U2493 (.IN1(n6988), .IN2(n2320), .IN3(\key_mem[2][122] ), .IN4(n6846), .Q(n3503)
          );
   AO22X1 U2494 (.IN1(n6869), .IN2(n2320), .IN3(\key_mem[3][122] ), .IN4(n6866), .Q(n3504)
          );
   AO22X1 U2495 (.IN1(n7288), .IN2(n2320), .IN3(\key_mem[4][122] ), .IN4(n6918), .Q(n3505)
          );
   AO22X1 U2496 (.IN1(n7274), .IN2(n2320), .IN3(\key_mem[5][122] ), .IN4(n7269), .Q(n3506)
          );
   AO22X1 U2497 (.IN1(n7266), .IN2(n2320), .IN3(\key_mem[6][122] ), .IN4(n7259), .Q(n3507)
          );
   AO22X1 U2498 (.IN1(n7014), .IN2(n2320), .IN3(\key_mem[7][122] ), .IN4(n7236), .Q(n3508)
          );
   AO22X1 U2499 (.IN1(n6752), .IN2(n2320), .IN3(\key_mem[8][122] ), .IN4(n6724), .Q(n3509)
          );
   AO22X1 U2500 (.IN1(n7218), .IN2(n2320), .IN3(\key_mem[9][122] ), .IN4(n7007), .Q(n3510)
          );
   AO22X1 U2501 (.IN1(n6799), .IN2(n2320), .IN3(\key_mem[10][122] ), .IN4(n6771), .Q(n3511)
          );
   AO22X1 U2502 (.IN1(n7194), .IN2(n2320), .IN3(\key_mem[11][122] ), .IN4(n7002), .Q(n3512)
          );
   AO22X1 U2503 (.IN1(n7186), .IN2(n2320), .IN3(\key_mem[12][122] ), .IN4(n6830), .Q(n3513)
          );
   AO22X1 U2504 (.IN1(n7173), .IN2(n2320), .IN3(\key_mem[13][122] ), .IN4(n6997), .Q(n3514)
          );
   AO22X1 U2505 (.IN1(n6996), .IN2(n2320), .IN3(\key_mem[14][122] ), .IN4(n7165), .Q(n3515)
          );
   AO221X1 U2506 (.IN1(n7126), .IN2(n2321), .IN3(key[250]), .IN4(n7292), .IN5(n2322), .Q(
          n2320));
   AO222X1 U2507 (.IN1(n7118), .IN2(n2323), .IN3(key[122]), .IN4(n7071), .IN5(n7038), .IN6(
          n2324), .Q(n2322));
   AO22X1 U2508 (.IN1(n7293), .IN2(n2325), .IN3(\key_mem[0][121] ), .IN4(n6938), .Q(n3516)
          );
   AO22X1 U2509 (.IN1(n6811), .IN2(n2325), .IN3(\key_mem[1][121] ), .IN4(n6821), .Q(n3517)
          );
   AO22X1 U2510 (.IN1(n6852), .IN2(n2325), .IN3(\key_mem[2][121] ), .IN4(n6843), .Q(n3518)
          );
   AO22X1 U2511 (.IN1(n6870), .IN2(n2325), .IN3(\key_mem[3][121] ), .IN4(n6877), .Q(n3519)
          );
   AO22X1 U2512 (.IN1(n6888), .IN2(n2325), .IN3(\key_mem[4][121] ), .IN4(n7021), .Q(n3520)
          );
   AO22X1 U2513 (.IN1(n7279), .IN2(n2325), .IN3(\key_mem[5][121] ), .IN4(n7269), .Q(n3521)
          );
   AO22X1 U2514 (.IN1(n7017), .IN2(n2325), .IN3(\key_mem[6][121] ), .IN4(n7254), .Q(n3522)
          );
   AO22X1 U2515 (.IN1(n7013), .IN2(n2325), .IN3(\key_mem[7][121] ), .IN4(n7237), .Q(n3523)
          );
   AO22X1 U2516 (.IN1(n6754), .IN2(n2325), .IN3(\key_mem[8][121] ), .IN4(n6747), .Q(n3524)
          );
   AO22X1 U2517 (.IN1(n7223), .IN2(n2325), .IN3(\key_mem[9][121] ), .IN4(n7212), .Q(n3525)
          );
   AO22X1 U2518 (.IN1(n6801), .IN2(n2325), .IN3(\key_mem[10][121] ), .IN4(n6794), .Q(n3526)
          );
   AO22X1 U2519 (.IN1(n7199), .IN2(n2325), .IN3(\key_mem[11][121] ), .IN4(n7188), .Q(n3527)
          );
   AO22X1 U2520 (.IN1(n6831), .IN2(n2325), .IN3(\key_mem[12][121] ), .IN4(n6834), .Q(n3528)
          );
   AO22X1 U2521 (.IN1(n7178), .IN2(n2325), .IN3(\key_mem[13][121] ), .IN4(n7167), .Q(n3529)
          );
   AO22X1 U2522 (.IN1(n6995), .IN2(n2325), .IN3(\key_mem[14][121] ), .IN4(n7157), .Q(n3530)
          );
   AO221X1 U2523 (.IN1(n7126), .IN2(n2326), .IN3(key[249]), .IN4(n7312), .IN5(n2327), .Q(
          n2325));
   AO222X1 U2524 (.IN1(n7117), .IN2(n2328), .IN3(key[121]), .IN4(n7071), .IN5(n7038), .IN6(
          n2329), .Q(n2327));
   AO22X1 U2525 (.IN1(n7306), .IN2(n2330), .IN3(\key_mem[0][120] ), .IN4(n6938), .Q(n3531)
          );
   AO22X1 U2526 (.IN1(n6927), .IN2(n2330), .IN3(\key_mem[1][120] ), .IN4(n6819), .Q(n3532)
          );
   AO22X1 U2527 (.IN1(n6988), .IN2(n2330), .IN3(\key_mem[2][120] ), .IN4(n6845), .Q(n3533)
          );
   AO22X1 U2528 (.IN1(n6870), .IN2(n2330), .IN3(\key_mem[3][120] ), .IN4(n6866), .Q(n3534)
          );
   AO22X1 U2529 (.IN1(n6886), .IN2(n2330), .IN3(\key_mem[4][120] ), .IN4(n7284), .Q(n3535)
          );
   AO22X1 U2530 (.IN1(n6974), .IN2(n2330), .IN3(\key_mem[5][120] ), .IN4(n7269), .Q(n3536)
          );
   AO22X1 U2531 (.IN1(n6969), .IN2(n2330), .IN3(\key_mem[6][120] ), .IN4(n7257), .Q(n3537)
          );
   AO22X1 U2532 (.IN1(n7246), .IN2(n2330), .IN3(\key_mem[7][120] ), .IN4(n7243), .Q(n3538)
          );
   AO22X1 U2533 (.IN1(n6750), .IN2(n2330), .IN3(\key_mem[8][120] ), .IN4(n6721), .Q(n3539)
          );
   AO22X1 U2534 (.IN1(n6976), .IN2(n2330), .IN3(\key_mem[9][120] ), .IN4(n7213), .Q(n3540)
          );
   AO22X1 U2535 (.IN1(n6797), .IN2(n2330), .IN3(\key_mem[10][120] ), .IN4(n6768), .Q(n3541)
          );
   AO22X1 U2536 (.IN1(n6978), .IN2(n2330), .IN3(\key_mem[11][120] ), .IN4(n7189), .Q(n3542)
          );
   AO22X1 U2537 (.IN1(n6827), .IN2(n2330), .IN3(\key_mem[12][120] ), .IN4(n7185), .Q(n3543)
          );
   AO22X1 U2538 (.IN1(n6980), .IN2(n2330), .IN3(\key_mem[13][120] ), .IN4(n7168), .Q(n3544)
          );
   AO22X1 U2539 (.IN1(n6992), .IN2(n2330), .IN3(\key_mem[14][120] ), .IN4(n7154), .Q(n3545)
          );
   AO221X1 U2540 (.IN1(n7126), .IN2(n2331), .IN3(key[248]), .IN4(n7301), .IN5(n2332), .Q(
          n2330));
   AO222X1 U2541 (.IN1(n7117), .IN2(n2333), .IN3(key[120]), .IN4(n7071), .IN5(n7038), .IN6(
          n2334), .Q(n2332));
   AO22X1 U2542 (.IN1(n7311), .IN2(n2335), .IN3(\key_mem[0][119] ), .IN4(n6937), .Q(n3546)
          );
   AO22X1 U2543 (.IN1(n6809), .IN2(n2335), .IN3(\key_mem[1][119] ), .IN4(n6820), .Q(n3547)
          );
   AO22X1 U2544 (.IN1(n6988), .IN2(n2335), .IN3(\key_mem[2][119] ), .IN4(n6845), .Q(n3548)
          );
   AO22X1 U2545 (.IN1(n6875), .IN2(n2335), .IN3(\key_mem[3][119] ), .IN4(n6863), .Q(n3549)
          );
   AO22X1 U2546 (.IN1(n6888), .IN2(n2335), .IN3(\key_mem[4][119] ), .IN4(n6917), .Q(n3550)
          );
   AO22X1 U2547 (.IN1(n7279), .IN2(n2335), .IN3(\key_mem[5][119] ), .IN4(n7270), .Q(n3551)
          );
   AO22X1 U2548 (.IN1(n7263), .IN2(n2335), .IN3(\key_mem[6][119] ), .IN4(n7255), .Q(n3552)
          );
   AO22X1 U2549 (.IN1(n7013), .IN2(n2335), .IN3(\key_mem[7][119] ), .IN4(n7238), .Q(n3553)
          );
   AO22X1 U2550 (.IN1(n6754), .IN2(n2335), .IN3(\key_mem[8][119] ), .IN4(n6738), .Q(n3554)
          );
   AO22X1 U2551 (.IN1(n7223), .IN2(n2335), .IN3(\key_mem[9][119] ), .IN4(n7216), .Q(n3555)
          );
   AO22X1 U2552 (.IN1(n6801), .IN2(n2335), .IN3(\key_mem[10][119] ), .IN4(n6785), .Q(n3556)
          );
   AO22X1 U2553 (.IN1(n7199), .IN2(n2335), .IN3(\key_mem[11][119] ), .IN4(n7192), .Q(n3557)
          );
   AO22X1 U2554 (.IN1(n6826), .IN2(n2335), .IN3(\key_mem[12][119] ), .IN4(n6833), .Q(n3558)
          );
   AO22X1 U2555 (.IN1(n7178), .IN2(n2335), .IN3(\key_mem[13][119] ), .IN4(n7171), .Q(n3559)
          );
   AO22X1 U2556 (.IN1(n7158), .IN2(n2335), .IN3(\key_mem[14][119] ), .IN4(n7155), .Q(n3560)
          );
   AO221X1 U2557 (.IN1(n7126), .IN2(n2336), .IN3(key[247]), .IN4(n7307), .IN5(n2337), .Q(
          n2335));
   AO222X1 U2558 (.IN1(n7117), .IN2(n2338), .IN3(key[119]), .IN4(n7071), .IN5(n7038), .IN6(
          n2339), .Q(n2337));
   AO22X1 U2559 (.IN1(n7309), .IN2(n2340), .IN3(\key_mem[0][118] ), .IN4(n6937), .Q(n3561)
          );
   AO22X1 U2561 (.IN1(n6988), .IN2(n2340), .IN3(\key_mem[2][118] ), .IN4(n6859), .Q(n3563)
          );
   AO22X1 U2562 (.IN1(n6875), .IN2(n2340), .IN3(\key_mem[3][118] ), .IN4(n6866), .Q(n3564)
          );
   AO22X1 U2563 (.IN1(n6916), .IN2(n2340), .IN3(\key_mem[4][118] ), .IN4(n7284), .Q(n3565)
          );
   AO22X1 U2564 (.IN1(n7280), .IN2(n2340), .IN3(\key_mem[5][118] ), .IN4(n7282), .Q(n3566)
          );
   AO22X1 U2565 (.IN1(n7264), .IN2(n2340), .IN3(\key_mem[6][118] ), .IN4(n7251), .Q(n3567)
          );
   AO22X1 U2566 (.IN1(n7013), .IN2(n2340), .IN3(\key_mem[7][118] ), .IN4(n7239), .Q(n3568)
          );
   AO22X1 U2567 (.IN1(n6750), .IN2(n2340), .IN3(\key_mem[8][118] ), .IN4(n6721), .Q(n3569)
          );
   AO22X1 U2568 (.IN1(n7224), .IN2(n2340), .IN3(\key_mem[9][118] ), .IN4(n7214), .Q(n3570)
          );
   AO22X1 U2569 (.IN1(n6797), .IN2(n2340), .IN3(\key_mem[10][118] ), .IN4(n6768), .Q(n3571)
          );
   AO22X1 U2570 (.IN1(n7200), .IN2(n2340), .IN3(\key_mem[11][118] ), .IN4(n7190), .Q(n3572)
          );
   AO22X1 U2571 (.IN1(n6987), .IN2(n2340), .IN3(\key_mem[12][118] ), .IN4(n7184), .Q(n3573)
          );
   AO22X1 U2572 (.IN1(n7179), .IN2(n2340), .IN3(\key_mem[13][118] ), .IN4(n7169), .Q(n3574)
          );
   AO22X1 U2573 (.IN1(n7159), .IN2(n2340), .IN3(\key_mem[14][118] ), .IN4(n7147), .Q(n3575)
          );
   AO222X1 U2575 (.IN1(n7117), .IN2(n2343), .IN3(key[118]), .IN4(n7071), .IN5(n7038), .IN6(
          n2344), .Q(n2342));
   AO22X1 U2576 (.IN1(n2276), .IN2(n2345), .IN3(\key_mem[0][117] ), .IN4(n6937), .Q(n3576)
          );
   AO22X1 U2577 (.IN1(n6812), .IN2(n2345), .IN3(\key_mem[1][117] ), .IN4(n6821), .Q(n3577)
          );
   AO22X1 U2578 (.IN1(n6852), .IN2(n2345), .IN3(\key_mem[2][117] ), .IN4(n6849), .Q(n3578)
          );
   AO22X1 U2579 (.IN1(n6875), .IN2(n2345), .IN3(\key_mem[3][117] ), .IN4(n6877), .Q(n3579)
          );
   AO22X1 U2580 (.IN1(n6916), .IN2(n2345), .IN3(\key_mem[4][117] ), .IN4(n6915), .Q(n3580)
          );
   AO22X1 U2581 (.IN1(n7274), .IN2(n2345), .IN3(\key_mem[5][117] ), .IN4(n7272), .Q(n3581)
          );
   AO22X1 U2582 (.IN1(n7266), .IN2(n2345), .IN3(\key_mem[6][117] ), .IN4(n2283), .Q(n3582)
          );
   AO22X1 U2583 (.IN1(n7245), .IN2(n2345), .IN3(\key_mem[7][117] ), .IN4(n7240), .Q(n3583)
          );
   AO22X1 U2584 (.IN1(n6751), .IN2(n2345), .IN3(\key_mem[8][117] ), .IN4(n6716), .Q(n3584)
          );
   AO22X1 U2585 (.IN1(n7218), .IN2(n2345), .IN3(\key_mem[9][117] ), .IN4(n7212), .Q(n3585)
          );
   AO22X1 U2586 (.IN1(n6798), .IN2(n2345), .IN3(\key_mem[10][117] ), .IN4(n6763), .Q(n3586)
          );
   AO22X1 U2587 (.IN1(n7194), .IN2(n2345), .IN3(\key_mem[11][117] ), .IN4(n7188), .Q(n3587)
          );
   AO22X1 U2588 (.IN1(n7183), .IN2(n2345), .IN3(\key_mem[12][117] ), .IN4(n6983), .Q(n3588)
          );
   AO22X1 U2589 (.IN1(n7173), .IN2(n2345), .IN3(\key_mem[13][117] ), .IN4(n7167), .Q(n3589)
          );
   AO22X1 U2590 (.IN1(n7164), .IN2(n2345), .IN3(\key_mem[14][117] ), .IN4(n7165), .Q(n3590)
          );
   AO221X1 U2591 (.IN1(n7126), .IN2(n2346), .IN3(key[245]), .IN4(n7303), .IN5(n2347), .Q(
          n2345));
   AO222X1 U2592 (.IN1(n7117), .IN2(n2348), .IN3(key[117]), .IN4(n7071), .IN5(n7038), .IN6(
          n2349), .Q(n2347));
   AO22X1 U2593 (.IN1(n7308), .IN2(n2350), .IN3(\key_mem[0][116] ), .IN4(n6937), .Q(n3591)
          );
   AO22X1 U2594 (.IN1(n6927), .IN2(n2350), .IN3(\key_mem[1][116] ), .IN4(n6821), .Q(n3592)
          );
   AO22X1 U2595 (.IN1(n6853), .IN2(n2350), .IN3(\key_mem[2][116] ), .IN4(n6851), .Q(n3593)
          );
   AO22X1 U2596 (.IN1(n6874), .IN2(n2350), .IN3(\key_mem[3][116] ), .IN4(n6861), .Q(n3594)
          );
   AO22X1 U2597 (.IN1(n7286), .IN2(n2350), .IN3(\key_mem[4][116] ), .IN4(n7021), .Q(n3595)
          );
   AO22X1 U2598 (.IN1(n7275), .IN2(n2350), .IN3(\key_mem[5][116] ), .IN4(n7018), .Q(n3596)
          );
   AO22X1 U2599 (.IN1(n7017), .IN2(n2350), .IN3(\key_mem[6][116] ), .IN4(n7015), .Q(n3597)
          );
   AO22X1 U2600 (.IN1(n7249), .IN2(n2350), .IN3(\key_mem[7][116] ), .IN4(n2284), .Q(n3598)
          );
   AO22X1 U2601 (.IN1(n6752), .IN2(n2350), .IN3(\key_mem[8][116] ), .IN4(n6737), .Q(n3599)
          );
   AO22X1 U2602 (.IN1(n7219), .IN2(n2350), .IN3(\key_mem[9][116] ), .IN4(n7216), .Q(n3600)
          );
   AO22X1 U2603 (.IN1(n6799), .IN2(n2350), .IN3(\key_mem[10][116] ), .IN4(n6784), .Q(n3601)
          );
   AO22X1 U2604 (.IN1(n7195), .IN2(n2350), .IN3(\key_mem[11][116] ), .IN4(n7192), .Q(n3602)
          );
   AO22X1 U2605 (.IN1(n6829), .IN2(n2350), .IN3(\key_mem[12][116] ), .IN4(n6830), .Q(n3603)
          );
   AO22X1 U2606 (.IN1(n7174), .IN2(n2350), .IN3(\key_mem[13][116] ), .IN4(n7171), .Q(n3604)
          );
   AO22X1 U2607 (.IN1(n6992), .IN2(n2350), .IN3(\key_mem[14][116] ), .IN4(n6994), .Q(n3605)
          );
   AO221X1 U2608 (.IN1(n7126), .IN2(n2351), .IN3(key[244]), .IN4(n7301), .IN5(n2352), .Q(
          n2350));
   AO222X1 U2609 (.IN1(n7117), .IN2(n2353), .IN3(key[116]), .IN4(n7071), .IN5(n7038), .IN6(
          n2354), .Q(n2352));
   AO22X1 U2610 (.IN1(n7293), .IN2(n2355), .IN3(\key_mem[0][115] ), .IN4(n6937), .Q(n3606)
          );
   AO22X1 U2611 (.IN1(n6811), .IN2(n2355), .IN3(\key_mem[1][115] ), .IN4(n6822), .Q(n3607)
          );
   AO22X1 U2612 (.IN1(n6852), .IN2(n2355), .IN3(\key_mem[2][115] ), .IN4(n6844), .Q(n3608)
          );
   AO22X1 U2613 (.IN1(n6874), .IN2(n2355), .IN3(\key_mem[3][115] ), .IN4(n6867), .Q(n3609)
          );
   AO22X1 U2614 (.IN1(n6921), .IN2(n2355), .IN3(\key_mem[4][115] ), .IN4(n6915), .Q(n3610)
          );
   AO22X1 U2615 (.IN1(n7275), .IN2(n2355), .IN3(\key_mem[5][115] ), .IN4(n7273), .Q(n3611)
          );
   AO22X1 U2616 (.IN1(n6969), .IN2(n2355), .IN3(\key_mem[6][115] ), .IN4(n2283), .Q(n3612)
          );
   AO22X1 U2617 (.IN1(n7250), .IN2(n2355), .IN3(\key_mem[7][115] ), .IN4(n2284), .Q(n3613)
          );
   AO22X1 U2618 (.IN1(n6751), .IN2(n2355), .IN3(\key_mem[8][115] ), .IN4(n6727), .Q(n3614)
          );
   AO22X1 U2619 (.IN1(n7219), .IN2(n2355), .IN3(\key_mem[9][115] ), .IN4(n7217), .Q(n3615)
          );
   AO22X1 U2620 (.IN1(n6798), .IN2(n2355), .IN3(\key_mem[10][115] ), .IN4(n6774), .Q(n3616)
          );
   AO22X1 U2621 (.IN1(n7195), .IN2(n2355), .IN3(\key_mem[11][115] ), .IN4(n7193), .Q(n3617)
          );
   AO22X1 U2622 (.IN1(n6987), .IN2(n2355), .IN3(\key_mem[12][115] ), .IN4(n6983), .Q(n3618)
          );
   AO22X1 U2623 (.IN1(n7174), .IN2(n2355), .IN3(\key_mem[13][115] ), .IN4(n7172), .Q(n3619)
          );
   AO22X1 U2624 (.IN1(n7163), .IN2(n2355), .IN3(\key_mem[14][115] ), .IN4(n7148), .Q(n3620)
          );
   AO221X1 U2625 (.IN1(n7127), .IN2(n2356), .IN3(key[243]), .IN4(n7300), .IN5(n2357), .Q(
          n2355));
   AO222X1 U2626 (.IN1(n7117), .IN2(n2358), .IN3(key[115]), .IN4(n7072), .IN5(n7039), .IN6(
          n2359), .Q(n2357));
   AO22X1 U2627 (.IN1(n7294), .IN2(n2360), .IN3(\key_mem[0][114] ), .IN4(n6937), .Q(n3621)
          );
   AO22X1 U2628 (.IN1(n6812), .IN2(n2360), .IN3(\key_mem[1][114] ), .IN4(n6823), .Q(n3622)
          );
   AO22X1 U2629 (.IN1(n6853), .IN2(n2360), .IN3(\key_mem[2][114] ), .IN4(n6846), .Q(n3623)
          );
   AO22X1 U2630 (.IN1(n6869), .IN2(n2360), .IN3(\key_mem[3][114] ), .IN4(n6864), .Q(n3624)
          );
   AO22X1 U2631 (.IN1(n6888), .IN2(n2360), .IN3(\key_mem[4][114] ), .IN4(n7289), .Q(n3625)
          );
   AO22X1 U2632 (.IN1(n7280), .IN2(n2360), .IN3(\key_mem[5][114] ), .IN4(n7273), .Q(n3626)
          );
   AO22X1 U2633 (.IN1(n7264), .IN2(n2360), .IN3(\key_mem[6][114] ), .IN4(n7015), .Q(n3627)
          );
   AO22X1 U2634 (.IN1(n7248), .IN2(n2360), .IN3(\key_mem[7][114] ), .IN4(n7238), .Q(n3628)
          );
   AO22X1 U2635 (.IN1(n6754), .IN2(n2360), .IN3(\key_mem[8][114] ), .IN4(n6735), .Q(n3629)
          );
   AO22X1 U2636 (.IN1(n7224), .IN2(n2360), .IN3(\key_mem[9][114] ), .IN4(n7213), .Q(n3630)
          );
   AO22X1 U2637 (.IN1(n6801), .IN2(n2360), .IN3(\key_mem[10][114] ), .IN4(n6782), .Q(n3631)
          );
   AO22X1 U2638 (.IN1(n7200), .IN2(n2360), .IN3(\key_mem[11][114] ), .IN4(n7189), .Q(n3632)
          );
   AO22X1 U2639 (.IN1(n6837), .IN2(n2360), .IN3(\key_mem[12][114] ), .IN4(n2289), .Q(n3633)
          );
   AO22X1 U2640 (.IN1(n7179), .IN2(n2360), .IN3(\key_mem[13][114] ), .IN4(n7168), .Q(n3634)
          );
   AO22X1 U2641 (.IN1(n7158), .IN2(n2360), .IN3(\key_mem[14][114] ), .IN4(n7147), .Q(n3635)
          );
   AO222X1 U2643 (.IN1(n7117), .IN2(n2363), .IN3(key[114]), .IN4(n7072), .IN5(n7039), .IN6(
          n2364), .Q(n2362));
   AO22X1 U2644 (.IN1(n7305), .IN2(n2365), .IN3(\key_mem[0][113] ), .IN4(n6937), .Q(n3636)
          );
   AO22X1 U2645 (.IN1(n6810), .IN2(n2365), .IN3(\key_mem[1][113] ), .IN4(n6819), .Q(n3637)
          );
   AO22X1 U2646 (.IN1(n6858), .IN2(n2365), .IN3(\key_mem[2][113] ), .IN4(n6851), .Q(n3638)
          );
   AO22X1 U2647 (.IN1(n6874), .IN2(n2365), .IN3(\key_mem[3][113] ), .IN4(n6867), .Q(n3639)
          );
   AO22X1 U2648 (.IN1(n6887), .IN2(n2365), .IN3(\key_mem[4][113] ), .IN4(n7021), .Q(n3640)
          );
   AO22X1 U2649 (.IN1(n7283), .IN2(n2365), .IN3(\key_mem[5][113] ), .IN4(n7271), .Q(n3641)
          );
   AO22X1 U2650 (.IN1(n7264), .IN2(n2365), .IN3(\key_mem[6][113] ), .IN4(n7258), .Q(n3642)
          );
   AO22X1 U2651 (.IN1(n7247), .IN2(n2365), .IN3(\key_mem[7][113] ), .IN4(n7241), .Q(n3643)
          );
   AO22X1 U2652 (.IN1(n6752), .IN2(n2365), .IN3(\key_mem[8][113] ), .IN4(n6726), .Q(n3644)
          );
   AO22X1 U2653 (.IN1(n7227), .IN2(n2365), .IN3(\key_mem[9][113] ), .IN4(n7214), .Q(n3645)
          );
   AO22X1 U2654 (.IN1(n6799), .IN2(n2365), .IN3(\key_mem[10][113] ), .IN4(n6773), .Q(n3646)
          );
   AO22X1 U2655 (.IN1(n7203), .IN2(n2365), .IN3(\key_mem[11][113] ), .IN4(n7190), .Q(n3647)
          );
   AO22X1 U2656 (.IN1(n6840), .IN2(n2365), .IN3(\key_mem[12][113] ), .IN4(n6981), .Q(n3648)
          );
   AO22X1 U2657 (.IN1(n7182), .IN2(n2365), .IN3(\key_mem[13][113] ), .IN4(n7169), .Q(n3649)
          );
   AO22X1 U2658 (.IN1(n7159), .IN2(n2365), .IN3(\key_mem[14][113] ), .IN4(n7153), .Q(n3650)
          );
   AO221X1 U2659 (.IN1(n7127), .IN2(n2366), .IN3(key[241]), .IN4(n7296), .IN5(n2367), .Q(
          n2365));
   AO222X1 U2660 (.IN1(n7117), .IN2(n2368), .IN3(key[113]), .IN4(n7072), .IN5(n7039), .IN6(
          n2369), .Q(n2367));
   AO22X1 U2661 (.IN1(n7290), .IN2(n2370), .IN3(\key_mem[0][112] ), .IN4(n6937), .Q(n3651)
          );
   AO22X1 U2662 (.IN1(n6927), .IN2(n2370), .IN3(\key_mem[1][112] ), .IN4(n6820), .Q(n3652)
          );
   AO22X1 U2663 (.IN1(n6852), .IN2(n2370), .IN3(\key_mem[2][112] ), .IN4(n6845), .Q(n3653)
          );
   AO22X1 U2664 (.IN1(n6875), .IN2(n2370), .IN3(\key_mem[3][112] ), .IN4(n6867), .Q(n3654)
          );
   AO22X1 U2665 (.IN1(n6921), .IN2(n2370), .IN3(\key_mem[4][112] ), .IN4(n6918), .Q(n3655)
          );
   AO22X1 U2666 (.IN1(n6974), .IN2(n2370), .IN3(\key_mem[5][112] ), .IN4(n7272), .Q(n3656)
          );
   AO22X1 U2667 (.IN1(n7264), .IN2(n2370), .IN3(\key_mem[6][112] ), .IN4(n7251), .Q(n3657)
          );
   AO22X1 U2668 (.IN1(n7246), .IN2(n2370), .IN3(\key_mem[7][112] ), .IN4(n7241), .Q(n3658)
          );
   AO22X1 U2669 (.IN1(n6754), .IN2(n2370), .IN3(\key_mem[8][112] ), .IN4(n6722), .Q(n3659)
          );
   AO22X1 U2670 (.IN1(n6976), .IN2(n2370), .IN3(\key_mem[9][112] ), .IN4(n7214), .Q(n3660)
          );
   AO22X1 U2671 (.IN1(n6801), .IN2(n2370), .IN3(\key_mem[10][112] ), .IN4(n6769), .Q(n3661)
          );
   AO22X1 U2672 (.IN1(n6978), .IN2(n2370), .IN3(\key_mem[11][112] ), .IN4(n7190), .Q(n3662)
          );
   AO22X1 U2673 (.IN1(n7001), .IN2(n2370), .IN3(\key_mem[12][112] ), .IN4(n6981), .Q(n3663)
          );
   AO22X1 U2674 (.IN1(n6980), .IN2(n2370), .IN3(\key_mem[13][112] ), .IN4(n7169), .Q(n3664)
          );
   AO22X1 U2675 (.IN1(n7162), .IN2(n2370), .IN3(\key_mem[14][112] ), .IN4(n7156), .Q(n3665)
          );
   AO221X1 U2676 (.IN1(n7127), .IN2(n2371), .IN3(key[240]), .IN4(n7299), .IN5(n2372), .Q(
          n2370));
   AO222X1 U2677 (.IN1(n7117), .IN2(n2373), .IN3(key[112]), .IN4(n7072), .IN5(n7039), .IN6(
          n2374), .Q(n2372));
   AO22X1 U2678 (.IN1(n7300), .IN2(n2375), .IN3(\key_mem[0][111] ), .IN4(n6937), .Q(n3666)
          );
   AO22X1 U2679 (.IN1(n6809), .IN2(n2375), .IN3(\key_mem[1][111] ), .IN4(n6821), .Q(n3667)
          );
   AO22X1 U2680 (.IN1(n6852), .IN2(n2375), .IN3(\key_mem[2][111] ), .IN4(n6851), .Q(n3668)
          );
   AO22X1 U2681 (.IN1(n6874), .IN2(n2375), .IN3(\key_mem[3][111] ), .IN4(n6860), .Q(n3669)
          );
   AO22X1 U2682 (.IN1(n6920), .IN2(n2375), .IN3(\key_mem[4][111] ), .IN4(n7289), .Q(n3670)
          );
   AO22X1 U2683 (.IN1(n7276), .IN2(n2375), .IN3(\key_mem[5][111] ), .IN4(n7267), .Q(n3671)
          );
   AO22X1 U2684 (.IN1(n7016), .IN2(n2375), .IN3(\key_mem[6][111] ), .IN4(n7259), .Q(n3672)
          );
   AO22X1 U2685 (.IN1(n7245), .IN2(n2375), .IN3(\key_mem[7][111] ), .IN4(n7242), .Q(n3673)
          );
   AO22X1 U2686 (.IN1(n6754), .IN2(n2375), .IN3(\key_mem[8][111] ), .IN4(n6717), .Q(n3674)
          );
   AO22X1 U2687 (.IN1(n7220), .IN2(n2375), .IN3(\key_mem[9][111] ), .IN4(n7214), .Q(n3675)
          );
   AO22X1 U2688 (.IN1(n6801), .IN2(n2375), .IN3(\key_mem[10][111] ), .IN4(n6764), .Q(n3676)
          );
   AO22X1 U2689 (.IN1(n7196), .IN2(n2375), .IN3(\key_mem[11][111] ), .IN4(n7190), .Q(n3677)
          );
   AO22X1 U2690 (.IN1(n6986), .IN2(n2375), .IN3(\key_mem[12][111] ), .IN4(n6983), .Q(n3678)
          );
   AO22X1 U2691 (.IN1(n7175), .IN2(n2375), .IN3(\key_mem[13][111] ), .IN4(n7169), .Q(n3679)
          );
   AO22X1 U2692 (.IN1(n6996), .IN2(n2375), .IN3(\key_mem[14][111] ), .IN4(n7151), .Q(n3680)
          );
   AO221X1 U2693 (.IN1(n7127), .IN2(n2376), .IN3(key[239]), .IN4(n7298), .IN5(n2377), .Q(
          n2375));
   AO222X1 U2694 (.IN1(n7117), .IN2(n2378), .IN3(key[111]), .IN4(n7072), .IN5(n7039), .IN6(
          n2379), .Q(n2377));
   AO22X1 U2695 (.IN1(n7302), .IN2(n2380), .IN3(\key_mem[0][110] ), .IN4(n6937), .Q(n3681)
          );
   AO22X1 U2696 (.IN1(n6808), .IN2(n2380), .IN3(\key_mem[1][110] ), .IN4(n6821), .Q(n3682)
          );
   AO22X1 U2697 (.IN1(n6858), .IN2(n2380), .IN3(\key_mem[2][110] ), .IN4(n6842), .Q(n3683)
          );
   AO22X1 U2698 (.IN1(n6874), .IN2(n2380), .IN3(\key_mem[3][110] ), .IN4(n6865), .Q(n3684)
          );
   AO22X1 U2699 (.IN1(n6920), .IN2(n2380), .IN3(\key_mem[4][110] ), .IN4(n6925), .Q(n3685)
          );
   AO22X1 U2700 (.IN1(n7275), .IN2(n2380), .IN3(\key_mem[5][110] ), .IN4(n7270), .Q(n3686)
          );
   AO22X1 U2701 (.IN1(n6969), .IN2(n2380), .IN3(\key_mem[6][110] ), .IN4(n7258), .Q(n3687)
          );
   AO22X1 U2702 (.IN1(n7249), .IN2(n2380), .IN3(\key_mem[7][110] ), .IN4(n7240), .Q(n3688)
          );
   AO22X1 U2703 (.IN1(n6755), .IN2(n2380), .IN3(\key_mem[8][110] ), .IN4(n6717), .Q(n3689)
          );
   AO22X1 U2704 (.IN1(n7219), .IN2(n2380), .IN3(\key_mem[9][110] ), .IN4(n7211), .Q(n3690)
          );
   AO22X1 U2705 (.IN1(n6802), .IN2(n2380), .IN3(\key_mem[10][110] ), .IN4(n6764), .Q(n3691)
          );
   AO22X1 U2706 (.IN1(n7195), .IN2(n2380), .IN3(\key_mem[11][110] ), .IN4(n7187), .Q(n3692)
          );
   AO22X1 U2707 (.IN1(n6986), .IN2(n2380), .IN3(\key_mem[12][110] ), .IN4(n2289), .Q(n3693)
          );
   AO22X1 U2708 (.IN1(n7174), .IN2(n2380), .IN3(\key_mem[13][110] ), .IN4(n7166), .Q(n3694)
          );
   AO22X1 U2709 (.IN1(n6971), .IN2(n2380), .IN3(\key_mem[14][110] ), .IN4(n7149), .Q(n3695)
          );
   AO221X1 U2710 (.IN1(n7127), .IN2(n2381), .IN3(key[238]), .IN4(n7299), .IN5(n2382), .Q(
          n2380));
   AO222X1 U2711 (.IN1(n7117), .IN2(n2383), .IN3(key[110]), .IN4(n7072), .IN5(n7039), .IN6(
          n2384), .Q(n2382));
   AO22X1 U2712 (.IN1(n7312), .IN2(n2385), .IN3(\key_mem[0][109] ), .IN4(n6937), .Q(n3696)
          );
   AO22X1 U2713 (.IN1(n6811), .IN2(n2385), .IN3(\key_mem[1][109] ), .IN4(n6814), .Q(n3697)
          );
   AO22X1 U2714 (.IN1(n6857), .IN2(n2385), .IN3(\key_mem[2][109] ), .IN4(n6846), .Q(n3698)
          );
   AO22X1 U2715 (.IN1(n6875), .IN2(n2385), .IN3(\key_mem[3][109] ), .IN4(n6867), .Q(n3699)
          );
   AO22X1 U2716 (.IN1(n7287), .IN2(n2385), .IN3(\key_mem[4][109] ), .IN4(n6919), .Q(n3700)
          );
   AO22X1 U2717 (.IN1(n7277), .IN2(n2385), .IN3(\key_mem[5][109] ), .IN4(n7273), .Q(n3701)
          );
   AO22X1 U2718 (.IN1(n6970), .IN2(n2385), .IN3(\key_mem[6][109] ), .IN4(n7256), .Q(n3702)
          );
   AO22X1 U2719 (.IN1(n7249), .IN2(n2385), .IN3(\key_mem[7][109] ), .IN4(n7242), .Q(n3703)
          );
   AO22X1 U2720 (.IN1(n6755), .IN2(n2385), .IN3(\key_mem[8][109] ), .IN4(n6725), .Q(n3704)
          );
   AO22X1 U2721 (.IN1(n7221), .IN2(n2385), .IN3(\key_mem[9][109] ), .IN4(n7007), .Q(n3705)
          );
   AO22X1 U2722 (.IN1(n6802), .IN2(n2385), .IN3(\key_mem[10][109] ), .IN4(n6772), .Q(n3706)
          );
   AO22X1 U2723 (.IN1(n7197), .IN2(n2385), .IN3(\key_mem[11][109] ), .IN4(n7002), .Q(n3707)
          );
   AO22X1 U2724 (.IN1(n6832), .IN2(n2385), .IN3(\key_mem[12][109] ), .IN4(n7000), .Q(n3708)
          );
   AO22X1 U2725 (.IN1(n7176), .IN2(n2385), .IN3(\key_mem[13][109] ), .IN4(n6997), .Q(n3709)
          );
   AO22X1 U2726 (.IN1(n6972), .IN2(n2385), .IN3(\key_mem[14][109] ), .IN4(n7165), .Q(n3710)
          );
   AO222X1 U2728 (.IN1(n7117), .IN2(n2388), .IN3(key[109]), .IN4(n7072), .IN5(n7039), .IN6(
          n2389), .Q(n2387));
   AO22X1 U2729 (.IN1(n7303), .IN2(n2390), .IN3(\key_mem[0][108] ), .IN4(n6937), .Q(n3711)
          );
   AO22X1 U2730 (.IN1(n6813), .IN2(n2390), .IN3(\key_mem[1][108] ), .IN4(n6817), .Q(n3712)
          );
   AO22X1 U2731 (.IN1(n6854), .IN2(n2390), .IN3(\key_mem[2][108] ), .IN4(n6842), .Q(n3713)
          );
   AO22X1 U2732 (.IN1(n6874), .IN2(n2390), .IN3(\key_mem[3][108] ), .IN4(n6876), .Q(n3714)
          );
   AO22X1 U2733 (.IN1(n6886), .IN2(n2390), .IN3(\key_mem[4][108] ), .IN4(n6914), .Q(n3715)
          );
   AO22X1 U2734 (.IN1(n7277), .IN2(n2390), .IN3(\key_mem[5][108] ), .IN4(n7273), .Q(n3716)
          );
   AO22X1 U2735 (.IN1(n7016), .IN2(n2390), .IN3(\key_mem[6][108] ), .IN4(n7255), .Q(n3717)
          );
   AO22X1 U2736 (.IN1(n7244), .IN2(n2390), .IN3(\key_mem[7][108] ), .IN4(n2284), .Q(n3718)
          );
   AO22X1 U2737 (.IN1(n6748), .IN2(n2390), .IN3(\key_mem[8][108] ), .IN4(n6718), .Q(n3719)
          );
   AO22X1 U2738 (.IN1(n7221), .IN2(n2390), .IN3(\key_mem[9][108] ), .IN4(n7217), .Q(n3720)
          );
   AO22X1 U2739 (.IN1(n6795), .IN2(n2390), .IN3(\key_mem[10][108] ), .IN4(n6765), .Q(n3721)
          );
   AO22X1 U2740 (.IN1(n7197), .IN2(n2390), .IN3(\key_mem[11][108] ), .IN4(n7193), .Q(n3722)
          );
   AO22X1 U2741 (.IN1(n6832), .IN2(n2390), .IN3(\key_mem[12][108] ), .IN4(n6828), .Q(n3723)
          );
   AO22X1 U2742 (.IN1(n7176), .IN2(n2390), .IN3(\key_mem[13][108] ), .IN4(n7172), .Q(n3724)
          );
   AO22X1 U2743 (.IN1(n7163), .IN2(n2390), .IN3(\key_mem[14][108] ), .IN4(n7150), .Q(n3725)
          );
   AO221X1 U2744 (.IN1(n7127), .IN2(n2391), .IN3(key[236]), .IN4(n7292), .IN5(n2392), .Q(
          n2390));
   AO222X1 U2745 (.IN1(n7116), .IN2(n2393), .IN3(key[108]), .IN4(n7072), .IN5(n7039), .IN6(
          n2394), .Q(n2392));
   AO22X1 U2746 (.IN1(n7301), .IN2(n2395), .IN3(\key_mem[0][107] ), .IN4(n6936), .Q(n3726)
          );
   AO22X1 U2747 (.IN1(n6812), .IN2(n2395), .IN3(\key_mem[1][107] ), .IN4(n6815), .Q(n3727)
          );
   AO22X1 U2748 (.IN1(n6855), .IN2(n2395), .IN3(\key_mem[2][107] ), .IN4(n6859), .Q(n3728)
          );
   AO22X1 U2749 (.IN1(n6871), .IN2(n2395), .IN3(\key_mem[3][107] ), .IN4(n6860), .Q(n3729)
          );
   AO22X1 U2750 (.IN1(n6887), .IN2(n2395), .IN3(\key_mem[4][107] ), .IN4(n6917), .Q(n3730)
          );
   AO22X1 U2751 (.IN1(n7280), .IN2(n2395), .IN3(\key_mem[5][107] ), .IN4(n7282), .Q(n3731)
          );
   AO22X1 U2752 (.IN1(n6969), .IN2(n2395), .IN3(\key_mem[6][107] ), .IN4(n7254), .Q(n3732)
          );
   AO22X1 U2753 (.IN1(n7245), .IN2(n2395), .IN3(\key_mem[7][107] ), .IN4(n7012), .Q(n3733)
          );
   AO22X1 U2754 (.IN1(n6755), .IN2(n2395), .IN3(\key_mem[8][107] ), .IN4(n6737), .Q(n3734)
          );
   AO22X1 U2755 (.IN1(n7224), .IN2(n2395), .IN3(\key_mem[9][107] ), .IN4(n7226), .Q(n3735)
          );
   AO22X1 U2756 (.IN1(n6802), .IN2(n2395), .IN3(\key_mem[10][107] ), .IN4(n6784), .Q(n3736)
          );
   AO22X1 U2757 (.IN1(n7200), .IN2(n2395), .IN3(\key_mem[11][107] ), .IN4(n7202), .Q(n3737)
          );
   AO22X1 U2758 (.IN1(n6827), .IN2(n2395), .IN3(\key_mem[12][107] ), .IN4(n6984), .Q(n3738)
          );
   AO22X1 U2759 (.IN1(n7179), .IN2(n2395), .IN3(\key_mem[13][107] ), .IN4(n7181), .Q(n3739)
          );
   AO22X1 U2760 (.IN1(n6996), .IN2(n2395), .IN3(\key_mem[14][107] ), .IN4(n6994), .Q(n3740)
          );
   AO222X1 U2762 (.IN1(n7116), .IN2(n2398), .IN3(key[107]), .IN4(n7072), .IN5(n7039), .IN6(
          n2399), .Q(n2397));
   AO22X1 U2763 (.IN1(n7308), .IN2(n2400), .IN3(\key_mem[0][106] ), .IN4(n6936), .Q(n3741)
          );
   AO22X1 U2764 (.IN1(n6811), .IN2(n2400), .IN3(\key_mem[1][106] ), .IN4(n6814), .Q(n3742)
          );
   AO22X1 U2765 (.IN1(n6853), .IN2(n2400), .IN3(\key_mem[2][106] ), .IN4(n6849), .Q(n3743)
          );
   AO22X1 U2766 (.IN1(n6871), .IN2(n2400), .IN3(\key_mem[3][106] ), .IN4(n6861), .Q(n3744)
          );
   AO22X1 U2767 (.IN1(n7288), .IN2(n2400), .IN3(\key_mem[4][106] ), .IN4(n6925), .Q(n3745)
          );
   AO22X1 U2768 (.IN1(n7278), .IN2(n2400), .IN3(\key_mem[5][106] ), .IN4(n7281), .Q(n3746)
          );
   AO22X1 U2769 (.IN1(n6970), .IN2(n2400), .IN3(\key_mem[6][106] ), .IN4(n7255), .Q(n3747)
          );
   AO22X1 U2770 (.IN1(n7244), .IN2(n2400), .IN3(\key_mem[7][106] ), .IN4(n7243), .Q(n3748)
          );
   AO22X1 U2771 (.IN1(n6752), .IN2(n2400), .IN3(\key_mem[8][106] ), .IN4(n6726), .Q(n3749)
          );
   AO22X1 U2772 (.IN1(n7222), .IN2(n2400), .IN3(\key_mem[9][106] ), .IN4(n7225), .Q(n3750)
          );
   AO22X1 U2773 (.IN1(n6799), .IN2(n2400), .IN3(\key_mem[10][106] ), .IN4(n6773), .Q(n3751)
          );
   AO22X1 U2774 (.IN1(n7198), .IN2(n2400), .IN3(\key_mem[11][106] ), .IN4(n7201), .Q(n3752)
          );
   AO22X1 U2775 (.IN1(n6986), .IN2(n2400), .IN3(\key_mem[12][106] ), .IN4(n7184), .Q(n3753)
          );
   AO22X1 U2776 (.IN1(n7177), .IN2(n2400), .IN3(\key_mem[13][106] ), .IN4(n7180), .Q(n3754)
          );
   AO22X1 U2777 (.IN1(n6995), .IN2(n2400), .IN3(\key_mem[14][106] ), .IN4(n7148), .Q(n3755)
          );
   AO222X1 U2779 (.IN1(n7116), .IN2(n2403), .IN3(key[106]), .IN4(n7072), .IN5(n7039), .IN6(
          n2404), .Q(n2402));
   AO22X1 U2780 (.IN1(n7309), .IN2(n2405), .IN3(\key_mem[0][105] ), .IN4(n6936), .Q(n3756)
          );
   AO22X1 U2781 (.IN1(n6927), .IN2(n2405), .IN3(\key_mem[1][105] ), .IN4(n6819), .Q(n3757)
          );
   AO22X1 U2782 (.IN1(n6855), .IN2(n2405), .IN3(\key_mem[2][105] ), .IN4(n6859), .Q(n3758)
          );
   AO22X1 U2783 (.IN1(n6872), .IN2(n2405), .IN3(\key_mem[3][105] ), .IN4(n6861), .Q(n3759)
          );
   AO22X1 U2784 (.IN1(n6990), .IN2(n2405), .IN3(\key_mem[4][105] ), .IN4(n7021), .Q(n3760)
          );
   AO22X1 U2785 (.IN1(n7019), .IN2(n2405), .IN3(\key_mem[5][105] ), .IN4(n7270), .Q(n3761)
          );
   AO22X1 U2786 (.IN1(n7265), .IN2(n2405), .IN3(\key_mem[6][105] ), .IN4(n7252), .Q(n3762)
          );
   AO22X1 U2787 (.IN1(n7014), .IN2(n2405), .IN3(\key_mem[7][105] ), .IN4(n7235), .Q(n3763)
          );
   AO22X1 U2788 (.IN1(n6758), .IN2(n2405), .IN3(\key_mem[8][105] ), .IN4(n6727), .Q(n3764)
          );
   AO22X1 U2789 (.IN1(n7008), .IN2(n2405), .IN3(\key_mem[9][105] ), .IN4(n7212), .Q(n3765)
          );
   AO22X1 U2790 (.IN1(n6805), .IN2(n2405), .IN3(\key_mem[10][105] ), .IN4(n6774), .Q(n3766)
          );
   AO22X1 U2791 (.IN1(n7003), .IN2(n2405), .IN3(\key_mem[11][105] ), .IN4(n7188), .Q(n3767)
          );
   AO22X1 U2792 (.IN1(n6835), .IN2(n2405), .IN3(\key_mem[12][105] ), .IN4(n6830), .Q(n3768)
          );
   AO22X1 U2793 (.IN1(n6998), .IN2(n2405), .IN3(\key_mem[13][105] ), .IN4(n7167), .Q(n3769)
          );
   AO22X1 U2794 (.IN1(n7160), .IN2(n2405), .IN3(\key_mem[14][105] ), .IN4(n7148), .Q(n3770)
          );
   AO222X1 U2796 (.IN1(n7116), .IN2(n2408), .IN3(key[105]), .IN4(n7072), .IN5(n7039), .IN6(
          n2409), .Q(n2407));
   AO22X1 U2797 (.IN1(n7307), .IN2(n2410), .IN3(\key_mem[0][104] ), .IN4(n6936), .Q(n3771)
          );
   AO22X1 U2798 (.IN1(n6809), .IN2(n2410), .IN3(\key_mem[1][104] ), .IN4(n6820), .Q(n3772)
          );
   AO22X1 U2799 (.IN1(n6857), .IN2(n2410), .IN3(\key_mem[2][104] ), .IN4(n6847), .Q(n3773)
          );
   AO22X1 U2800 (.IN1(n6871), .IN2(n2410), .IN3(\key_mem[3][104] ), .IN4(n6860), .Q(n3774)
          );
   AO22X1 U2801 (.IN1(n6889), .IN2(n2410), .IN3(\key_mem[4][104] ), .IN4(n6890), .Q(n3775)
          );
   AO22X1 U2802 (.IN1(n7280), .IN2(n2410), .IN3(\key_mem[5][104] ), .IN4(n7273), .Q(n3776)
          );
   AO22X1 U2803 (.IN1(n6970), .IN2(n2410), .IN3(\key_mem[6][104] ), .IN4(n7253), .Q(n3777)
          );
   AO22X1 U2804 (.IN1(n7013), .IN2(n2410), .IN3(\key_mem[7][104] ), .IN4(n7236), .Q(n3778)
          );
   AO22X1 U2805 (.IN1(n6756), .IN2(n2410), .IN3(\key_mem[8][104] ), .IN4(n6735), .Q(n3779)
          );
   AO22X1 U2806 (.IN1(n7224), .IN2(n2410), .IN3(\key_mem[9][104] ), .IN4(n7212), .Q(n3780)
          );
   AO22X1 U2807 (.IN1(n6803), .IN2(n2410), .IN3(\key_mem[10][104] ), .IN4(n6782), .Q(n3781)
          );
   AO22X1 U2808 (.IN1(n7200), .IN2(n2410), .IN3(\key_mem[11][104] ), .IN4(n7188), .Q(n3782)
          );
   AO22X1 U2809 (.IN1(n6826), .IN2(n2410), .IN3(\key_mem[12][104] ), .IN4(n7185), .Q(n3783)
          );
   AO22X1 U2810 (.IN1(n7179), .IN2(n2410), .IN3(\key_mem[13][104] ), .IN4(n7167), .Q(n3784)
          );
   AO22X1 U2811 (.IN1(n6971), .IN2(n2410), .IN3(\key_mem[14][104] ), .IN4(n7154), .Q(n3785)
          );
   AO222X1 U2813 (.IN1(n7116), .IN2(n2413), .IN3(key[104]), .IN4(n7072), .IN5(n7039), .IN6(
          n2414), .Q(n2412));
   AO22X1 U2814 (.IN1(n7302), .IN2(n2415), .IN3(\key_mem[0][103] ), .IN4(n6936), .Q(n3786)
          );
   AO22X1 U2815 (.IN1(n6808), .IN2(n2415), .IN3(\key_mem[1][103] ), .IN4(n6815), .Q(n3787)
          );
   AO22X1 U2816 (.IN1(n6854), .IN2(n2415), .IN3(\key_mem[2][103] ), .IN4(n6849), .Q(n3788)
          );
   AO22X1 U2817 (.IN1(n6870), .IN2(n2415), .IN3(\key_mem[3][103] ), .IN4(n6866), .Q(n3789)
          );
   AO22X1 U2818 (.IN1(n7022), .IN2(n2415), .IN3(\key_mem[4][103] ), .IN4(n6914), .Q(n3790)
          );
   AO22X1 U2819 (.IN1(n7278), .IN2(n2415), .IN3(\key_mem[5][103] ), .IN4(n7271), .Q(n3791)
          );
   AO22X1 U2820 (.IN1(n7266), .IN2(n2415), .IN3(\key_mem[6][103] ), .IN4(n7256), .Q(n3792)
          );
   AO22X1 U2821 (.IN1(n7249), .IN2(n2415), .IN3(\key_mem[7][103] ), .IN4(n7012), .Q(n3793)
          );
   AO22X1 U2822 (.IN1(n6755), .IN2(n2415), .IN3(\key_mem[8][103] ), .IN4(n6722), .Q(n3794)
          );
   AO22X1 U2823 (.IN1(n7222), .IN2(n2415), .IN3(\key_mem[9][103] ), .IN4(n7215), .Q(n3795)
          );
   AO22X1 U2824 (.IN1(n6802), .IN2(n2415), .IN3(\key_mem[10][103] ), .IN4(n6769), .Q(n3796)
          );
   AO22X1 U2825 (.IN1(n7198), .IN2(n2415), .IN3(\key_mem[11][103] ), .IN4(n7191), .Q(n3797)
          );
   AO22X1 U2826 (.IN1(n6829), .IN2(n2415), .IN3(\key_mem[12][103] ), .IN4(n7184), .Q(n3798)
          );
   AO22X1 U2827 (.IN1(n7177), .IN2(n2415), .IN3(\key_mem[13][103] ), .IN4(n7170), .Q(n3799)
          );
   AO22X1 U2828 (.IN1(n7164), .IN2(n2415), .IN3(\key_mem[14][103] ), .IN4(n7155), .Q(n3800)
          );
   AO221X1 U2829 (.IN1(n7128), .IN2(n2416), .IN3(key[231]), .IN4(n7292), .IN5(n2417), .Q(
          n2415));
   AO222X1 U2830 (.IN1(n7116), .IN2(n2418), .IN3(key[103]), .IN4(n7073), .IN5(n7040), .IN6(
          n2419), .Q(n2417));
   AO22X1 U2831 (.IN1(n7302), .IN2(n2420), .IN3(\key_mem[0][102] ), .IN4(n6936), .Q(n3801)
          );
   AO22X1 U2832 (.IN1(n6810), .IN2(n2420), .IN3(\key_mem[1][102] ), .IN4(n6816), .Q(n3802)
          );
   AO22X1 U2833 (.IN1(n6853), .IN2(n2420), .IN3(\key_mem[2][102] ), .IN4(n6851), .Q(n3803)
          );
   AO22X1 U2834 (.IN1(n6871), .IN2(n2420), .IN3(\key_mem[3][102] ), .IN4(n6861), .Q(n3804)
          );
   AO22X1 U2835 (.IN1(n7288), .IN2(n2420), .IN3(\key_mem[4][102] ), .IN4(n6914), .Q(n3805)
          );
   AO22X1 U2836 (.IN1(n7020), .IN2(n2420), .IN3(\key_mem[5][102] ), .IN4(n7282), .Q(n3806)
          );
   AO22X1 U2837 (.IN1(n7266), .IN2(n2420), .IN3(\key_mem[6][102] ), .IN4(n7258), .Q(n3807)
          );
   AO22X1 U2838 (.IN1(n7244), .IN2(n2420), .IN3(\key_mem[7][102] ), .IN4(n7012), .Q(n3808)
          );
   AO22X1 U2839 (.IN1(n6756), .IN2(n2420), .IN3(\key_mem[8][102] ), .IN4(n6721), .Q(n3809)
          );
   AO22X1 U2840 (.IN1(n7009), .IN2(n2420), .IN3(\key_mem[9][102] ), .IN4(n7226), .Q(n3810)
          );
   AO22X1 U2841 (.IN1(n6803), .IN2(n2420), .IN3(\key_mem[10][102] ), .IN4(n6768), .Q(n3811)
          );
   AO22X1 U2842 (.IN1(n7004), .IN2(n2420), .IN3(\key_mem[11][102] ), .IN4(n7202), .Q(n3812)
          );
   AO22X1 U2843 (.IN1(n6837), .IN2(n2420), .IN3(\key_mem[12][102] ), .IN4(n7185), .Q(n3813)
          );
   AO22X1 U2844 (.IN1(n6999), .IN2(n2420), .IN3(\key_mem[13][102] ), .IN4(n7181), .Q(n3814)
          );
   AO22X1 U2845 (.IN1(n6995), .IN2(n2420), .IN3(\key_mem[14][102] ), .IN4(n7147), .Q(n3815)
          );
   AO221X1 U2846 (.IN1(n7128), .IN2(n2421), .IN3(key[230]), .IN4(n2276), .IN5(n2422), .Q(
          n2420));
   AO222X1 U2847 (.IN1(n7116), .IN2(n2423), .IN3(key[102]), .IN4(n7073), .IN5(n7040), .IN6(
          n2424), .Q(n2422));
   AO22X1 U2848 (.IN1(n7301), .IN2(n2425), .IN3(\key_mem[0][101] ), .IN4(n6936), .Q(n3816)
          );
   AO22X1 U2849 (.IN1(n6809), .IN2(n2425), .IN3(\key_mem[1][101] ), .IN4(n6815), .Q(n3817)
          );
   AO22X1 U2850 (.IN1(n6853), .IN2(n2425), .IN3(\key_mem[2][101] ), .IN4(n6843), .Q(n3818)
          );
   AO22X1 U2851 (.IN1(n6871), .IN2(n2425), .IN3(\key_mem[3][101] ), .IN4(n6868), .Q(n3819)
          );
   AO22X1 U2852 (.IN1(n6916), .IN2(n2425), .IN3(\key_mem[4][101] ), .IN4(n6918), .Q(n3820)
          );
   AO22X1 U2853 (.IN1(n6973), .IN2(n2425), .IN3(\key_mem[5][101] ), .IN4(n7270), .Q(n3821)
          );
   AO22X1 U2854 (.IN1(n7266), .IN2(n2425), .IN3(\key_mem[6][101] ), .IN4(n7257), .Q(n3822)
          );
   AO22X1 U2855 (.IN1(n7250), .IN2(n2425), .IN3(\key_mem[7][101] ), .IN4(n7239), .Q(n3823)
          );
   AO22X1 U2856 (.IN1(n6757), .IN2(n2425), .IN3(\key_mem[8][101] ), .IN4(n6727), .Q(n3824)
          );
   AO22X1 U2857 (.IN1(n6975), .IN2(n2425), .IN3(\key_mem[9][101] ), .IN4(n7211), .Q(n3825)
          );
   AO22X1 U2858 (.IN1(n6804), .IN2(n2425), .IN3(\key_mem[10][101] ), .IN4(n6774), .Q(n3826)
          );
   AO22X1 U2859 (.IN1(n6977), .IN2(n2425), .IN3(\key_mem[11][101] ), .IN4(n7187), .Q(n3827)
          );
   AO22X1 U2860 (.IN1(n6829), .IN2(n2425), .IN3(\key_mem[12][101] ), .IN4(n6985), .Q(n3828)
          );
   AO22X1 U2861 (.IN1(n6979), .IN2(n2425), .IN3(\key_mem[13][101] ), .IN4(n7166), .Q(n3829)
          );
   AO22X1 U2862 (.IN1(n6992), .IN2(n2425), .IN3(\key_mem[14][101] ), .IN4(n7165), .Q(n3830)
          );
   AO221X1 U2863 (.IN1(n7128), .IN2(n2426), .IN3(key[229]), .IN4(n7309), .IN5(n2427), .Q(
          n2425));
   AO222X1 U2864 (.IN1(n7116), .IN2(n2428), .IN3(key[101]), .IN4(n7073), .IN5(n7040), .IN6(
          n2429), .Q(n2427));
   AO22X1 U2865 (.IN1(n7300), .IN2(n2430), .IN3(\key_mem[0][100] ), .IN4(n6936), .Q(n3831)
          );
   AO22X1 U2866 (.IN1(n6813), .IN2(n2430), .IN3(\key_mem[1][100] ), .IN4(n6814), .Q(n3832)
          );
   AO22X1 U2867 (.IN1(n6855), .IN2(n2430), .IN3(\key_mem[2][100] ), .IN4(n6846), .Q(n3833)
          );
   AO22X1 U2868 (.IN1(n6872), .IN2(n2430), .IN3(\key_mem[3][100] ), .IN4(n6867), .Q(n3834)
          );
   AO22X1 U2869 (.IN1(n6921), .IN2(n2430), .IN3(\key_mem[4][100] ), .IN4(n7289), .Q(n3835)
          );
   AO22X1 U2870 (.IN1(n7279), .IN2(n2430), .IN3(\key_mem[5][100] ), .IN4(n7282), .Q(n3836)
          );
   AO22X1 U2871 (.IN1(n6970), .IN2(n2430), .IN3(\key_mem[6][100] ), .IN4(n7252), .Q(n3837)
          );
   AO22X1 U2872 (.IN1(n7250), .IN2(n2430), .IN3(\key_mem[7][100] ), .IN4(n7242), .Q(n3838)
          );
   AO22X1 U2873 (.IN1(n6758), .IN2(n2430), .IN3(\key_mem[8][100] ), .IN4(n6717), .Q(n3839)
          );
   AO22X1 U2874 (.IN1(n7223), .IN2(n2430), .IN3(\key_mem[9][100] ), .IN4(n7226), .Q(n3840)
          );
   AO22X1 U2875 (.IN1(n6805), .IN2(n2430), .IN3(\key_mem[10][100] ), .IN4(n6764), .Q(n3841)
          );
   AO22X1 U2876 (.IN1(n7199), .IN2(n2430), .IN3(\key_mem[11][100] ), .IN4(n7202), .Q(n3842)
          );
   AO22X1 U2877 (.IN1(n7186), .IN2(n2430), .IN3(\key_mem[12][100] ), .IN4(n7184), .Q(n3843)
          );
   AO22X1 U2878 (.IN1(n7178), .IN2(n2430), .IN3(\key_mem[13][100] ), .IN4(n7181), .Q(n3844)
          );
   AO22X1 U2879 (.IN1(n7158), .IN2(n2430), .IN3(\key_mem[14][100] ), .IN4(n6994), .Q(n3845)
          );
   AO221X1 U2880 (.IN1(n7128), .IN2(n2431), .IN3(key[228]), .IN4(n7312), .IN5(n2432), .Q(
          n2430));
   AO222X1 U2881 (.IN1(n7116), .IN2(n2433), .IN3(key[100]), .IN4(n7073), .IN5(n7040), .IN6(
          n2434), .Q(n2432));
   AO22X1 U2882 (.IN1(n7307), .IN2(n2435), .IN3(\key_mem[0][99] ), .IN4(n6936), .Q(n3846)
          );
   AO22X1 U2883 (.IN1(n6808), .IN2(n2435), .IN3(\key_mem[1][99] ), .IN4(n6825), .Q(n3847)
          );
   AO22X1 U2884 (.IN1(n6856), .IN2(n2435), .IN3(\key_mem[2][99] ), .IN4(n6851), .Q(n3848)
          );
   AO22X1 U2885 (.IN1(n6871), .IN2(n2435), .IN3(\key_mem[3][99] ), .IN4(n6866), .Q(n3849)
          );
   AO22X1 U2886 (.IN1(n7287), .IN2(n2435), .IN3(\key_mem[4][99] ), .IN4(n6925), .Q(n3850)
          );
   AO22X1 U2887 (.IN1(n7274), .IN2(n2435), .IN3(\key_mem[5][99] ), .IN4(n7281), .Q(n3851)
          );
   AO22X1 U2888 (.IN1(n7265), .IN2(n2435), .IN3(\key_mem[6][99] ), .IN4(n7255), .Q(n3852)
          );
   AO22X1 U2889 (.IN1(n7014), .IN2(n2435), .IN3(\key_mem[7][99] ), .IN4(n7237), .Q(n3853)
          );
   AO22X1 U2890 (.IN1(n6752), .IN2(n2435), .IN3(\key_mem[8][99] ), .IN4(n6721), .Q(n3854)
          );
   AO22X1 U2891 (.IN1(n7218), .IN2(n2435), .IN3(\key_mem[9][99] ), .IN4(n7225), .Q(n3855)
          );
   AO22X1 U2892 (.IN1(n6799), .IN2(n2435), .IN3(\key_mem[10][99] ), .IN4(n6768), .Q(n3856)
          );
   AO22X1 U2893 (.IN1(n7194), .IN2(n2435), .IN3(\key_mem[11][99] ), .IN4(n7201), .Q(n3857)
          );
   AO22X1 U2894 (.IN1(n6837), .IN2(n2435), .IN3(\key_mem[12][99] ), .IN4(n6984), .Q(n3858)
          );
   AO22X1 U2895 (.IN1(n7173), .IN2(n2435), .IN3(\key_mem[13][99] ), .IN4(n7180), .Q(n3859)
          );
   AO22X1 U2896 (.IN1(n6971), .IN2(n2435), .IN3(\key_mem[14][99] ), .IN4(n7148), .Q(n3860)
          );
   AO221X1 U2897 (.IN1(n7128), .IN2(n2436), .IN3(key[227]), .IN4(n7309), .IN5(n2437), .Q(
          n2435));
   AO222X1 U2898 (.IN1(n7116), .IN2(n2438), .IN3(key[99]), .IN4(n7073), .IN5(n7040), .IN6(
          n2439), .Q(n2437));
   AO22X1 U2899 (.IN1(n7306), .IN2(n2440), .IN3(\key_mem[0][98] ), .IN4(n6936), .Q(n3861)
          );
   AO22X1 U2900 (.IN1(n6809), .IN2(n2440), .IN3(\key_mem[1][98] ), .IN4(n6815), .Q(n3862)
          );
   AO22X1 U2901 (.IN1(n6988), .IN2(n2440), .IN3(\key_mem[2][98] ), .IN4(n6848), .Q(n3863)
          );
   AO22X1 U2902 (.IN1(n6872), .IN2(n2440), .IN3(\key_mem[3][98] ), .IN4(n6868), .Q(n3864)
          );
   AO22X1 U2903 (.IN1(n6924), .IN2(n2440), .IN3(\key_mem[4][98] ), .IN4(n7285), .Q(n3865)
          );
   AO22X1 U2904 (.IN1(n7280), .IN2(n2440), .IN3(\key_mem[5][98] ), .IN4(n7018), .Q(n3866)
          );
   AO22X1 U2905 (.IN1(n7265), .IN2(n2440), .IN3(\key_mem[6][98] ), .IN4(n7252), .Q(n3867)
          );
   AO22X1 U2906 (.IN1(n7250), .IN2(n2440), .IN3(\key_mem[7][98] ), .IN4(n7238), .Q(n3868)
          );
   AO22X1 U2907 (.IN1(n6757), .IN2(n2440), .IN3(\key_mem[8][98] ), .IN4(n6721), .Q(n3869)
          );
   AO22X1 U2908 (.IN1(n7224), .IN2(n2440), .IN3(\key_mem[9][98] ), .IN4(n7007), .Q(n3870)
          );
   AO22X1 U2909 (.IN1(n6804), .IN2(n2440), .IN3(\key_mem[10][98] ), .IN4(n6768), .Q(n3871)
          );
   AO22X1 U2910 (.IN1(n7200), .IN2(n2440), .IN3(\key_mem[11][98] ), .IN4(n7002), .Q(n3872)
          );
   AO22X1 U2911 (.IN1(n7186), .IN2(n2440), .IN3(\key_mem[12][98] ), .IN4(n6834), .Q(n3873)
          );
   AO22X1 U2912 (.IN1(n7179), .IN2(n2440), .IN3(\key_mem[13][98] ), .IN4(n6997), .Q(n3874)
          );
   AO22X1 U2913 (.IN1(n7164), .IN2(n2440), .IN3(\key_mem[14][98] ), .IN4(n7150), .Q(n3875)
          );
   AO221X1 U2914 (.IN1(n7128), .IN2(n2441), .IN3(key[226]), .IN4(n7307), .IN5(n2442), .Q(
          n2440));
   AO222X1 U2915 (.IN1(n7116), .IN2(n2443), .IN3(key[98]), .IN4(n7073), .IN5(n7040), .IN6(
          n2444), .Q(n2442));
   AO22X1 U2916 (.IN1(n7305), .IN2(n2445), .IN3(\key_mem[0][97] ), .IN4(n6936), .Q(n3876)
          );
   AO22X1 U2917 (.IN1(n6808), .IN2(n2445), .IN3(\key_mem[1][97] ), .IN4(n6825), .Q(n3877)
          );
   AO22X1 U2918 (.IN1(n6855), .IN2(n2445), .IN3(\key_mem[2][97] ), .IN4(n6842), .Q(n3878)
          );
   AO22X1 U2919 (.IN1(n6807), .IN2(n2445), .IN3(\key_mem[3][97] ), .IN4(n6865), .Q(n3879)
          );
   AO22X1 U2920 (.IN1(n7287), .IN2(n2445), .IN3(\key_mem[4][97] ), .IN4(n6917), .Q(n3880)
          );
   AO22X1 U2921 (.IN1(n7276), .IN2(n2445), .IN3(\key_mem[5][97] ), .IN4(n7268), .Q(n3881)
          );
   AO22X1 U2922 (.IN1(n7260), .IN2(n2445), .IN3(\key_mem[6][97] ), .IN4(n7254), .Q(n3882)
          );
   AO22X1 U2923 (.IN1(n7248), .IN2(n2445), .IN3(\key_mem[7][97] ), .IN4(n7239), .Q(n3883)
          );
   AO22X1 U2924 (.IN1(n6756), .IN2(n2445), .IN3(\key_mem[8][97] ), .IN4(n6725), .Q(n3884)
          );
   AO22X1 U2925 (.IN1(n7220), .IN2(n2445), .IN3(\key_mem[9][97] ), .IN4(n7212), .Q(n3885)
          );
   AO22X1 U2926 (.IN1(n6803), .IN2(n2445), .IN3(\key_mem[10][97] ), .IN4(n6772), .Q(n3886)
          );
   AO22X1 U2927 (.IN1(n7196), .IN2(n2445), .IN3(\key_mem[11][97] ), .IN4(n7188), .Q(n3887)
          );
   AO22X1 U2928 (.IN1(n7186), .IN2(n2445), .IN3(\key_mem[12][97] ), .IN4(n6981), .Q(n3888)
          );
   AO22X1 U2929 (.IN1(n7175), .IN2(n2445), .IN3(\key_mem[13][97] ), .IN4(n7167), .Q(n3889)
          );
   AO22X1 U2930 (.IN1(n7160), .IN2(n2445), .IN3(\key_mem[14][97] ), .IN4(n7151), .Q(n3890)
          );
   AO222X1 U2932 (.IN1(n7116), .IN2(n2448), .IN3(key[97]), .IN4(n7073), .IN5(n7040), .IN6(
          n2449), .Q(n2447));
   AO22X1 U2933 (.IN1(n2276), .IN2(n2450), .IN3(\key_mem[0][96] ), .IN4(n6936), .Q(n3891)
          );
   AO22X1 U2934 (.IN1(n6926), .IN2(n2450), .IN3(\key_mem[1][96] ), .IN4(n6814), .Q(n3892)
          );
   AO22X1 U2935 (.IN1(n6855), .IN2(n2450), .IN3(\key_mem[2][96] ), .IN4(n6845), .Q(n3893)
          );
   AO22X1 U2936 (.IN1(n6873), .IN2(n2450), .IN3(\key_mem[3][96] ), .IN4(n6865), .Q(n3894)
          );
   AO22X1 U2937 (.IN1(n6921), .IN2(n2450), .IN3(\key_mem[4][96] ), .IN4(n6890), .Q(n3895)
          );
   AO22X1 U2938 (.IN1(n7276), .IN2(n2450), .IN3(\key_mem[5][96] ), .IN4(n7272), .Q(n3896)
          );
   AO22X1 U2939 (.IN1(n7261), .IN2(n2450), .IN3(\key_mem[6][96] ), .IN4(n2283), .Q(n3897)
          );
   AO22X1 U2940 (.IN1(n7247), .IN2(n2450), .IN3(\key_mem[7][96] ), .IN4(n7240), .Q(n3898)
          );
   AO22X1 U2941 (.IN1(n6757), .IN2(n2450), .IN3(\key_mem[8][96] ), .IN4(n6724), .Q(n3899)
          );
   AO22X1 U2942 (.IN1(n7220), .IN2(n2450), .IN3(\key_mem[9][96] ), .IN4(n7215), .Q(n3900)
          );
   AO22X1 U2943 (.IN1(n6804), .IN2(n2450), .IN3(\key_mem[10][96] ), .IN4(n6771), .Q(n3901)
          );
   AO22X1 U2944 (.IN1(n7196), .IN2(n2450), .IN3(\key_mem[11][96] ), .IN4(n7191), .Q(n3902)
          );
   AO22X1 U2945 (.IN1(n6986), .IN2(n2450), .IN3(\key_mem[12][96] ), .IN4(n6841), .Q(n3903)
          );
   AO22X1 U2946 (.IN1(n7175), .IN2(n2450), .IN3(\key_mem[13][96] ), .IN4(n7170), .Q(n3904)
          );
   AO22X1 U2947 (.IN1(n7161), .IN2(n2450), .IN3(\key_mem[14][96] ), .IN4(n7148), .Q(n3905)
          );
   AO222X1 U2949 (.IN1(n7116), .IN2(n2453), .IN3(key[96]), .IN4(n7073), .IN5(n7040), .IN6(
          n2454), .Q(n2452));
   AO22X1 U2950 (.IN1(n7312), .IN2(n2455), .IN3(\key_mem[0][95] ), .IN4(n6935), .Q(n3906)
          );
   AO22X1 U2951 (.IN1(n6812), .IN2(n2455), .IN3(\key_mem[1][95] ), .IN4(n6816), .Q(n3907)
          );
   AO22X1 U2952 (.IN1(n6856), .IN2(n2455), .IN3(\key_mem[2][95] ), .IN4(n6849), .Q(n3908)
          );
   AO22X1 U2953 (.IN1(n6806), .IN2(n2455), .IN3(\key_mem[3][95] ), .IN4(n6861), .Q(n3909)
          );
   AO22X1 U2954 (.IN1(n6886), .IN2(n2455), .IN3(\key_mem[4][95] ), .IN4(n6914), .Q(n3910)
          );
   AO22X1 U2955 (.IN1(n7274), .IN2(n2455), .IN3(\key_mem[5][95] ), .IN4(n2282), .Q(n3911)
          );
   AO22X1 U2956 (.IN1(n7262), .IN2(n2455), .IN3(\key_mem[6][95] ), .IN4(n7015), .Q(n3912)
          );
   AO22X1 U2957 (.IN1(n7246), .IN2(n2455), .IN3(\key_mem[7][95] ), .IN4(n7241), .Q(n3913)
          );
   AO22X1 U2958 (.IN1(n6755), .IN2(n2455), .IN3(\key_mem[8][95] ), .IN4(n6741), .Q(n3914)
          );
   AO22X1 U2959 (.IN1(n7218), .IN2(n2455), .IN3(\key_mem[9][95] ), .IN4(n2286), .Q(n3915)
          );
   AO22X1 U2960 (.IN1(n6802), .IN2(n2455), .IN3(\key_mem[10][95] ), .IN4(n6788), .Q(n3916)
          );
   AO22X1 U2961 (.IN1(n7194), .IN2(n2455), .IN3(\key_mem[11][95] ), .IN4(n2288), .Q(n3917)
          );
   AO22X1 U2962 (.IN1(n6829), .IN2(n2455), .IN3(\key_mem[12][95] ), .IN4(n6841), .Q(n3918)
          );
   AO22X1 U2963 (.IN1(n7173), .IN2(n2455), .IN3(\key_mem[13][95] ), .IN4(n2290), .Q(n3919)
          );
   AO22X1 U2964 (.IN1(n6992), .IN2(n2455), .IN3(\key_mem[14][95] ), .IN4(n7149), .Q(n3920)
          );
   AO221X1 U2965 (.IN1(n7128), .IN2(n2456), .IN3(key[223]), .IN4(n7308), .IN5(n2457), .Q(
          n2455));
   AO222X1 U2966 (.IN1(n7115), .IN2(n2458), .IN3(key[95]), .IN4(n7073), .IN5(n7040), .IN6(
          n2459), .Q(n2457));
   AO22X1 U2967 (.IN1(n7305), .IN2(n2460), .IN3(\key_mem[0][94] ), .IN4(n6935), .Q(n3921)
          );
   AO22X1 U2968 (.IN1(n6809), .IN2(n2460), .IN3(\key_mem[1][94] ), .IN4(n6823), .Q(n3922)
          );
   AO22X1 U2969 (.IN1(n6858), .IN2(n2460), .IN3(\key_mem[2][94] ), .IN4(n6848), .Q(n3923)
          );
   AO22X1 U2970 (.IN1(n6872), .IN2(n2460), .IN3(\key_mem[3][94] ), .IN4(n6860), .Q(n3924)
          );
   AO22X1 U2971 (.IN1(n6887), .IN2(n2460), .IN3(\key_mem[4][94] ), .IN4(n6917), .Q(n3925)
          );
   AO22X1 U2972 (.IN1(n7020), .IN2(n2460), .IN3(\key_mem[5][94] ), .IN4(n7282), .Q(n3926)
          );
   AO22X1 U2973 (.IN1(n7263), .IN2(n2460), .IN3(\key_mem[6][94] ), .IN4(n7251), .Q(n3927)
          );
   AO22X1 U2974 (.IN1(n7245), .IN2(n2460), .IN3(\key_mem[7][94] ), .IN4(n7242), .Q(n3928)
          );
   AO22X1 U2975 (.IN1(n6756), .IN2(n2460), .IN3(\key_mem[8][94] ), .IN4(n6739), .Q(n3929)
          );
   AO22X1 U2976 (.IN1(n7009), .IN2(n2460), .IN3(\key_mem[9][94] ), .IN4(n7226), .Q(n3930)
          );
   AO22X1 U2977 (.IN1(n6803), .IN2(n2460), .IN3(\key_mem[10][94] ), .IN4(n6786), .Q(n3931)
          );
   AO22X1 U2978 (.IN1(n7004), .IN2(n2460), .IN3(\key_mem[11][94] ), .IN4(n7202), .Q(n3932)
          );
   AO22X1 U2979 (.IN1(n6987), .IN2(n2460), .IN3(\key_mem[12][94] ), .IN4(n6981), .Q(n3933)
          );
   AO22X1 U2980 (.IN1(n6999), .IN2(n2460), .IN3(\key_mem[13][94] ), .IN4(n7181), .Q(n3934)
          );
   AO22X1 U2981 (.IN1(n6971), .IN2(n2460), .IN3(\key_mem[14][94] ), .IN4(n7151), .Q(n3935)
          );
   AO221X1 U2982 (.IN1(n7128), .IN2(n2461), .IN3(key[222]), .IN4(n7302), .IN5(n2462), .Q(
          n2460));
   AO222X1 U2983 (.IN1(n7115), .IN2(n2463), .IN3(key[94]), .IN4(n7073), .IN5(n7040), .IN6(
          n2464), .Q(n2462));
   AO22X1 U2984 (.IN1(n7309), .IN2(n2465), .IN3(\key_mem[0][93] ), .IN4(n6935), .Q(n3936)
          );
   AO22X1 U2985 (.IN1(n6809), .IN2(n2465), .IN3(\key_mem[1][93] ), .IN4(n6814), .Q(n3937)
          );
   AO22X1 U2986 (.IN1(n6858), .IN2(n2465), .IN3(\key_mem[2][93] ), .IN4(n6846), .Q(n3938)
          );
   AO22X1 U2987 (.IN1(n6875), .IN2(n2465), .IN3(\key_mem[3][93] ), .IN4(n6861), .Q(n3939)
          );
   AO22X1 U2988 (.IN1(n6888), .IN2(n2465), .IN3(\key_mem[4][93] ), .IN4(n6917), .Q(n3940)
          );
   AO22X1 U2989 (.IN1(n7278), .IN2(n2465), .IN3(\key_mem[5][93] ), .IN4(n7281), .Q(n3941)
          );
   AO22X1 U2990 (.IN1(n7265), .IN2(n2465), .IN3(\key_mem[6][93] ), .IN4(n7251), .Q(n3942)
          );
   AO22X1 U2991 (.IN1(n7014), .IN2(n2465), .IN3(\key_mem[7][93] ), .IN4(n7236), .Q(n3943)
          );
   AO22X1 U2992 (.IN1(n6751), .IN2(n2465), .IN3(\key_mem[8][93] ), .IN4(n6730), .Q(n3944)
          );
   AO22X1 U2993 (.IN1(n7222), .IN2(n2465), .IN3(\key_mem[9][93] ), .IN4(n7225), .Q(n3945)
          );
   AO22X1 U2994 (.IN1(n6798), .IN2(n2465), .IN3(\key_mem[10][93] ), .IN4(n6777), .Q(n3946)
          );
   AO22X1 U2995 (.IN1(n7198), .IN2(n2465), .IN3(\key_mem[11][93] ), .IN4(n7201), .Q(n3947)
          );
   AO22X1 U2996 (.IN1(n6827), .IN2(n2465), .IN3(\key_mem[12][93] ), .IN4(n6985), .Q(n3948)
          );
   AO22X1 U2997 (.IN1(n7177), .IN2(n2465), .IN3(\key_mem[13][93] ), .IN4(n7180), .Q(n3949)
          );
   AO22X1 U2998 (.IN1(n7161), .IN2(n2465), .IN3(\key_mem[14][93] ), .IN4(n7155), .Q(n3950)
          );
   AO221X1 U2999 (.IN1(n7128), .IN2(n2466), .IN3(key[221]), .IN4(n7295), .IN5(n2467), .Q(
          n2465));
   AO222X1 U3000 (.IN1(n7115), .IN2(n2468), .IN3(key[93]), .IN4(n7073), .IN5(n7040), .IN6(
          n2469), .Q(n2467));
   AO22X1 U3001 (.IN1(n7311), .IN2(n2470), .IN3(\key_mem[0][92] ), .IN4(n6935), .Q(n3951)
          );
   AO22X1 U3002 (.IN1(n6811), .IN2(n2470), .IN3(\key_mem[1][92] ), .IN4(n6816), .Q(n3952)
          );
   AO22X1 U3003 (.IN1(n6852), .IN2(n2470), .IN3(\key_mem[2][92] ), .IN4(n6842), .Q(n3953)
          );
   AO22X1 U3004 (.IN1(n6872), .IN2(n2470), .IN3(\key_mem[3][92] ), .IN4(n6876), .Q(n3954)
          );
   AO22X1 U3005 (.IN1(n7288), .IN2(n2470), .IN3(\key_mem[4][92] ), .IN4(n6923), .Q(n3955)
          );
   AO22X1 U3006 (.IN1(n7020), .IN2(n2470), .IN3(\key_mem[5][92] ), .IN4(n7018), .Q(n3956)
          );
   AO22X1 U3007 (.IN1(n7017), .IN2(n2470), .IN3(\key_mem[6][92] ), .IN4(n7259), .Q(n3957)
          );
   AO22X1 U3008 (.IN1(n7248), .IN2(n2470), .IN3(\key_mem[7][92] ), .IN4(n7239), .Q(n3958)
          );
   AO22X1 U3009 (.IN1(n6750), .IN2(n2470), .IN3(\key_mem[8][92] ), .IN4(n6724), .Q(n3959)
          );
   AO22X1 U3010 (.IN1(n7009), .IN2(n2470), .IN3(\key_mem[9][92] ), .IN4(n7007), .Q(n3960)
          );
   AO22X1 U3011 (.IN1(n6797), .IN2(n2470), .IN3(\key_mem[10][92] ), .IN4(n6771), .Q(n3961)
          );
   AO22X1 U3012 (.IN1(n7004), .IN2(n2470), .IN3(\key_mem[11][92] ), .IN4(n7002), .Q(n3962)
          );
   AO22X1 U3013 (.IN1(n6831), .IN2(n2470), .IN3(\key_mem[12][92] ), .IN4(n7185), .Q(n3963)
          );
   AO22X1 U3014 (.IN1(n6999), .IN2(n2470), .IN3(\key_mem[13][92] ), .IN4(n6997), .Q(n3964)
          );
   AO22X1 U3015 (.IN1(n6972), .IN2(n2470), .IN3(\key_mem[14][92] ), .IN4(n7152), .Q(n3965)
          );
   AO221X1 U3016 (.IN1(n7128), .IN2(n2471), .IN3(key[220]), .IN4(n7303), .IN5(n2472), .Q(
          n2470));
   AO222X1 U3017 (.IN1(n7115), .IN2(n2473), .IN3(key[92]), .IN4(n7073), .IN5(n7040), .IN6(
          n2474), .Q(n2472));
   AO22X1 U3018 (.IN1(n7294), .IN2(n2475), .IN3(\key_mem[0][91] ), .IN4(n6935), .Q(n3966)
          );
   AO22X1 U3019 (.IN1(n6926), .IN2(n2475), .IN3(\key_mem[1][91] ), .IN4(n6817), .Q(n3967)
          );
   AO22X1 U3020 (.IN1(n6853), .IN2(n2475), .IN3(\key_mem[2][91] ), .IN4(n6843), .Q(n3968)
          );
   AO22X1 U3021 (.IN1(n6873), .IN2(n2475), .IN3(\key_mem[3][91] ), .IN4(n6877), .Q(n3969)
          );
   AO22X1 U3022 (.IN1(n7287), .IN2(n2475), .IN3(\key_mem[4][91] ), .IN4(n6914), .Q(n3970)
          );
   AO22X1 U3023 (.IN1(n7019), .IN2(n2475), .IN3(\key_mem[5][91] ), .IN4(n7269), .Q(n3971)
          );
   AO22X1 U3024 (.IN1(n7017), .IN2(n2475), .IN3(\key_mem[6][91] ), .IN4(n7258), .Q(n3972)
          );
   AO22X1 U3025 (.IN1(n7248), .IN2(n2475), .IN3(\key_mem[7][91] ), .IN4(n2284), .Q(n3973)
          );
   AO22X1 U3026 (.IN1(n6751), .IN2(n2475), .IN3(\key_mem[8][91] ), .IN4(n6730), .Q(n3974)
          );
   AO22X1 U3027 (.IN1(n7008), .IN2(n2475), .IN3(\key_mem[9][91] ), .IN4(n7212), .Q(n3975)
          );
   AO22X1 U3028 (.IN1(n6798), .IN2(n2475), .IN3(\key_mem[10][91] ), .IN4(n6777), .Q(n3976)
          );
   AO22X1 U3029 (.IN1(n7003), .IN2(n2475), .IN3(\key_mem[11][91] ), .IN4(n7188), .Q(n3977)
          );
   AO22X1 U3030 (.IN1(n6832), .IN2(n2475), .IN3(\key_mem[12][91] ), .IN4(n6828), .Q(n3978)
          );
   AO22X1 U3031 (.IN1(n6998), .IN2(n2475), .IN3(\key_mem[13][91] ), .IN4(n7167), .Q(n3979)
          );
   AO22X1 U3032 (.IN1(n7160), .IN2(n2475), .IN3(\key_mem[14][91] ), .IN4(n7149), .Q(n3980)
          );
   AO221X1 U3033 (.IN1(n7129), .IN2(n2476), .IN3(key[219]), .IN4(n7296), .IN5(n2477), .Q(
          n2475));
   AO222X1 U3034 (.IN1(n7115), .IN2(n2478), .IN3(key[91]), .IN4(n7074), .IN5(n7041), .IN6(
          n2479), .Q(n2477));
   AO22X1 U3035 (.IN1(n7291), .IN2(n2480), .IN3(\key_mem[0][90] ), .IN4(n6935), .Q(n3981)
          );
   AO22X1 U3036 (.IN1(n6813), .IN2(n2480), .IN3(\key_mem[1][90] ), .IN4(n6818), .Q(n3982)
          );
   AO22X1 U3037 (.IN1(n6858), .IN2(n2480), .IN3(\key_mem[2][90] ), .IN4(n6859), .Q(n3983)
          );
   AO22X1 U3038 (.IN1(n6806), .IN2(n2480), .IN3(\key_mem[3][90] ), .IN4(n6862), .Q(n3984)
          );
   AO22X1 U3039 (.IN1(n7288), .IN2(n2480), .IN3(\key_mem[4][90] ), .IN4(n7285), .Q(n3985)
          );
   AO22X1 U3040 (.IN1(n7283), .IN2(n2480), .IN3(\key_mem[5][90] ), .IN4(n7268), .Q(n3986)
          );
   AO22X1 U3041 (.IN1(n7017), .IN2(n2480), .IN3(\key_mem[6][90] ), .IN4(n7257), .Q(n3987)
          );
   AO22X1 U3042 (.IN1(n7013), .IN2(n2480), .IN3(\key_mem[7][90] ), .IN4(n7243), .Q(n3988)
          );
   AO22X1 U3043 (.IN1(n6752), .IN2(n2480), .IN3(\key_mem[8][90] ), .IN4(n6717), .Q(n3989)
          );
   AO22X1 U3044 (.IN1(n7227), .IN2(n2480), .IN3(\key_mem[9][90] ), .IN4(n7213), .Q(n3990)
          );
   AO22X1 U3045 (.IN1(n6799), .IN2(n2480), .IN3(\key_mem[10][90] ), .IN4(n6764), .Q(n3991)
          );
   AO22X1 U3046 (.IN1(n7203), .IN2(n2480), .IN3(\key_mem[11][90] ), .IN4(n7189), .Q(n3992)
          );
   AO22X1 U3047 (.IN1(n6827), .IN2(n2480), .IN3(\key_mem[12][90] ), .IN4(n7185), .Q(n3993)
          );
   AO22X1 U3048 (.IN1(n7182), .IN2(n2480), .IN3(\key_mem[13][90] ), .IN4(n7168), .Q(n3994)
          );
   AO22X1 U3049 (.IN1(n6972), .IN2(n2480), .IN3(\key_mem[14][90] ), .IN4(n7152), .Q(n3995)
          );
   AO221X1 U3050 (.IN1(n7129), .IN2(n2481), .IN3(key[218]), .IN4(n7299), .IN5(n2482), .Q(
          n2480));
   AO222X1 U3051 (.IN1(n7115), .IN2(n2483), .IN3(key[90]), .IN4(n7074), .IN5(n7041), .IN6(
          n2484), .Q(n2482));
   AO22X1 U3052 (.IN1(n7293), .IN2(n2485), .IN3(\key_mem[0][89] ), .IN4(n6935), .Q(n3996)
          );
   AO22X1 U3053 (.IN1(n6813), .IN2(n2485), .IN3(\key_mem[1][89] ), .IN4(n6815), .Q(n3997)
          );
   AO22X1 U3054 (.IN1(n6858), .IN2(n2485), .IN3(\key_mem[2][89] ), .IN4(n6848), .Q(n3998)
          );
   AO22X1 U3055 (.IN1(n6873), .IN2(n2485), .IN3(\key_mem[3][89] ), .IN4(n6862), .Q(n3999)
          );
   AO22X1 U3056 (.IN1(n6889), .IN2(n2485), .IN3(\key_mem[4][89] ), .IN4(n6915), .Q(n4000)
          );
   AO22X1 U3057 (.IN1(n6974), .IN2(n2485), .IN3(\key_mem[5][89] ), .IN4(n7268), .Q(n4001)
          );
   AO22X1 U3058 (.IN1(n7260), .IN2(n2485), .IN3(\key_mem[6][89] ), .IN4(n7256), .Q(n4002)
          );
   AO22X1 U3059 (.IN1(n7244), .IN2(n2485), .IN3(\key_mem[7][89] ), .IN4(n7243), .Q(n4003)
          );
   AO22X1 U3060 (.IN1(n6754), .IN2(n2485), .IN3(\key_mem[8][89] ), .IN4(n6719), .Q(n4004)
          );
   AO22X1 U3061 (.IN1(n6976), .IN2(n2485), .IN3(\key_mem[9][89] ), .IN4(n7213), .Q(n4005)
          );
   AO22X1 U3062 (.IN1(n6801), .IN2(n2485), .IN3(\key_mem[10][89] ), .IN4(n6766), .Q(n4006)
          );
   AO22X1 U3063 (.IN1(n6978), .IN2(n2485), .IN3(\key_mem[11][89] ), .IN4(n7189), .Q(n4007)
          );
   AO22X1 U3064 (.IN1(n6987), .IN2(n2485), .IN3(\key_mem[12][89] ), .IN4(n6828), .Q(n4008)
          );
   AO22X1 U3065 (.IN1(n6980), .IN2(n2485), .IN3(\key_mem[13][89] ), .IN4(n7168), .Q(n4009)
          );
   AO22X1 U3066 (.IN1(n7163), .IN2(n2485), .IN3(\key_mem[14][89] ), .IN4(n7153), .Q(n4010)
          );
   AO221X1 U3067 (.IN1(n7129), .IN2(n2486), .IN3(key[217]), .IN4(n7298), .IN5(n2487), .Q(
          n2485));
   AO222X1 U3068 (.IN1(n7115), .IN2(n2488), .IN3(key[89]), .IN4(n7074), .IN5(n7041), .IN6(
          n2489), .Q(n2487));
   AO22X1 U3069 (.IN1(n7294), .IN2(n2490), .IN3(\key_mem[0][88] ), .IN4(n6935), .Q(n4011)
          );
   AO22X1 U3070 (.IN1(n6927), .IN2(n2490), .IN3(\key_mem[1][88] ), .IN4(n6816), .Q(n4012)
          );
   AO22X1 U3071 (.IN1(n6988), .IN2(n2490), .IN3(\key_mem[2][88] ), .IN4(n6843), .Q(n4013)
          );
   AO22X1 U3072 (.IN1(n6806), .IN2(n2490), .IN3(\key_mem[3][88] ), .IN4(n6861), .Q(n4014)
          );
   AO22X1 U3073 (.IN1(n6916), .IN2(n2490), .IN3(\key_mem[4][88] ), .IN4(n6925), .Q(n4015)
          );
   AO22X1 U3074 (.IN1(n7277), .IN2(n2490), .IN3(\key_mem[5][88] ), .IN4(n7272), .Q(n4016)
          );
   AO22X1 U3075 (.IN1(n7261), .IN2(n2490), .IN3(\key_mem[6][88] ), .IN4(n7254), .Q(n4017)
          );
   AO22X1 U3076 (.IN1(n7014), .IN2(n2490), .IN3(\key_mem[7][88] ), .IN4(n7240), .Q(n4018)
          );
   AO22X1 U3077 (.IN1(n6757), .IN2(n2490), .IN3(\key_mem[8][88] ), .IN4(n6738), .Q(n4019)
          );
   AO22X1 U3078 (.IN1(n7221), .IN2(n2490), .IN3(\key_mem[9][88] ), .IN4(n7216), .Q(n4020)
          );
   AO22X1 U3079 (.IN1(n6804), .IN2(n2490), .IN3(\key_mem[10][88] ), .IN4(n6785), .Q(n4021)
          );
   AO22X1 U3080 (.IN1(n7197), .IN2(n2490), .IN3(\key_mem[11][88] ), .IN4(n7192), .Q(n4022)
          );
   AO22X1 U3081 (.IN1(n7183), .IN2(n2490), .IN3(\key_mem[12][88] ), .IN4(n7185), .Q(n4023)
          );
   AO22X1 U3082 (.IN1(n7176), .IN2(n2490), .IN3(\key_mem[13][88] ), .IN4(n7171), .Q(n4024)
          );
   AO22X1 U3083 (.IN1(n7159), .IN2(n2490), .IN3(\key_mem[14][88] ), .IN4(n7150), .Q(n4025)
          );
   AO221X1 U3084 (.IN1(n7129), .IN2(n2491), .IN3(key[216]), .IN4(n7297), .IN5(n2492), .Q(
          n2490));
   AO222X1 U3085 (.IN1(n7115), .IN2(n2493), .IN3(key[88]), .IN4(n7074), .IN5(n7041), .IN6(
          n2494), .Q(n2492));
   AO22X1 U3086 (.IN1(n7291), .IN2(n2495), .IN3(\key_mem[0][87] ), .IN4(n6935), .Q(n4026)
          );
   AO22X1 U3087 (.IN1(n6810), .IN2(n2495), .IN3(\key_mem[1][87] ), .IN4(n6818), .Q(n4027)
          );
   AO22X1 U3088 (.IN1(n6852), .IN2(n2495), .IN3(\key_mem[2][87] ), .IN4(n6844), .Q(n4028)
          );
   AO22X1 U3089 (.IN1(n6871), .IN2(n2495), .IN3(\key_mem[3][87] ), .IN4(n6866), .Q(n4029)
          );
   AO22X1 U3090 (.IN1(n6921), .IN2(n2495), .IN3(\key_mem[4][87] ), .IN4(n6925), .Q(n4030)
          );
   AO22X1 U3091 (.IN1(n7275), .IN2(n2495), .IN3(\key_mem[5][87] ), .IN4(n7281), .Q(n4031)
          );
   AO22X1 U3092 (.IN1(n7260), .IN2(n2495), .IN3(\key_mem[6][87] ), .IN4(n7253), .Q(n4032)
          );
   AO22X1 U3093 (.IN1(n7013), .IN2(n2495), .IN3(\key_mem[7][87] ), .IN4(n7235), .Q(n4033)
          );
   AO22X1 U3094 (.IN1(n6752), .IN2(n2495), .IN3(\key_mem[8][87] ), .IN4(n6729), .Q(n4034)
          );
   AO22X1 U3095 (.IN1(n7219), .IN2(n2495), .IN3(\key_mem[9][87] ), .IN4(n7225), .Q(n4035)
          );
   AO22X1 U3096 (.IN1(n6799), .IN2(n2495), .IN3(\key_mem[10][87] ), .IN4(n6776), .Q(n4036)
          );
   AO22X1 U3097 (.IN1(n7195), .IN2(n2495), .IN3(\key_mem[11][87] ), .IN4(n7201), .Q(n4037)
          );
   AO22X1 U3098 (.IN1(n6829), .IN2(n2495), .IN3(\key_mem[12][87] ), .IN4(n7184), .Q(n4038)
          );
   AO22X1 U3099 (.IN1(n7174), .IN2(n2495), .IN3(\key_mem[13][87] ), .IN4(n7180), .Q(n4039)
          );
   AO22X1 U3100 (.IN1(n7164), .IN2(n2495), .IN3(\key_mem[14][87] ), .IN4(n7151), .Q(n4040)
          );
   AO221X1 U3101 (.IN1(n7129), .IN2(n2496), .IN3(key[215]), .IN4(n7290), .IN5(n2497), .Q(
          n2495));
   AO222X1 U3102 (.IN1(n7115), .IN2(n2498), .IN3(key[87]), .IN4(n7074), .IN5(n7041), .IN6(
          n2499), .Q(n2497));
   AO22X1 U3103 (.IN1(n7298), .IN2(n2500), .IN3(\key_mem[0][86] ), .IN4(n6935), .Q(n4041)
          );
   AO22X1 U3104 (.IN1(n6813), .IN2(n2500), .IN3(\key_mem[1][86] ), .IN4(n6823), .Q(n4042)
          );
   AO22X1 U3105 (.IN1(n6857), .IN2(n2500), .IN3(\key_mem[2][86] ), .IN4(n6859), .Q(n4043)
          );
   AO22X1 U3106 (.IN1(n6807), .IN2(n2500), .IN3(\key_mem[3][86] ), .IN4(n6866), .Q(n4044)
          );
   AO22X1 U3107 (.IN1(n6924), .IN2(n2500), .IN3(\key_mem[4][86] ), .IN4(n6914), .Q(n4045)
          );
   AO22X1 U3108 (.IN1(n7278), .IN2(n2500), .IN3(\key_mem[5][86] ), .IN4(n7271), .Q(n4046)
          );
   AO22X1 U3109 (.IN1(n7264), .IN2(n2500), .IN3(\key_mem[6][86] ), .IN4(n7253), .Q(n4047)
          );
   AO22X1 U3110 (.IN1(n7249), .IN2(n2500), .IN3(\key_mem[7][86] ), .IN4(n7012), .Q(n4048)
          );
   AO22X1 U3111 (.IN1(n6757), .IN2(n2500), .IN3(\key_mem[8][86] ), .IN4(n6727), .Q(n4049)
          );
   AO22X1 U3112 (.IN1(n7222), .IN2(n2500), .IN3(\key_mem[9][86] ), .IN4(n7217), .Q(n4050)
          );
   AO22X1 U3113 (.IN1(n6804), .IN2(n2500), .IN3(\key_mem[10][86] ), .IN4(n6774), .Q(n4051)
          );
   AO22X1 U3114 (.IN1(n7198), .IN2(n2500), .IN3(\key_mem[11][86] ), .IN4(n7193), .Q(n4052)
          );
   AO22X1 U3115 (.IN1(n6827), .IN2(n2500), .IN3(\key_mem[12][86] ), .IN4(n6983), .Q(n4053)
          );
   AO22X1 U3116 (.IN1(n7177), .IN2(n2500), .IN3(\key_mem[13][86] ), .IN4(n7172), .Q(n4054)
          );
   AO22X1 U3117 (.IN1(n7162), .IN2(n2500), .IN3(\key_mem[14][86] ), .IN4(n7148), .Q(n4055)
          );
   AO221X1 U3118 (.IN1(n7129), .IN2(n2501), .IN3(key[214]), .IN4(n7293), .IN5(n2502), .Q(
          n2500));
   AO222X1 U3119 (.IN1(n7115), .IN2(n2503), .IN3(key[86]), .IN4(n7074), .IN5(n7041), .IN6(
          n2504), .Q(n2502));
   AO22X1 U3120 (.IN1(n7296), .IN2(n2505), .IN3(\key_mem[0][85] ), .IN4(n6935), .Q(n4056)
          );
   AO22X1 U3121 (.IN1(n6927), .IN2(n2505), .IN3(\key_mem[1][85] ), .IN4(n6824), .Q(n4057)
          );
   AO22X1 U3122 (.IN1(n6857), .IN2(n2505), .IN3(\key_mem[2][85] ), .IN4(n6848), .Q(n4058)
          );
   AO22X1 U3123 (.IN1(n6989), .IN2(n2505), .IN3(\key_mem[3][85] ), .IN4(n6864), .Q(n4059)
          );
   AO22X1 U3124 (.IN1(n7287), .IN2(n2505), .IN3(\key_mem[4][85] ), .IN4(n7285), .Q(n4060)
          );
   AO22X1 U3125 (.IN1(n7274), .IN2(n2505), .IN3(\key_mem[5][85] ), .IN4(n7268), .Q(n4061)
          );
   AO22X1 U3126 (.IN1(n7266), .IN2(n2505), .IN3(\key_mem[6][85] ), .IN4(n7257), .Q(n4062)
          );
   AO22X1 U3127 (.IN1(n7250), .IN2(n2505), .IN3(\key_mem[7][85] ), .IN4(n7243), .Q(n4063)
          );
   AO22X1 U3128 (.IN1(n6758), .IN2(n2505), .IN3(\key_mem[8][85] ), .IN4(n6729), .Q(n4064)
          );
   AO22X1 U3129 (.IN1(n7218), .IN2(n2505), .IN3(\key_mem[9][85] ), .IN4(n7213), .Q(n4065)
          );
   AO22X1 U3130 (.IN1(n6805), .IN2(n2505), .IN3(\key_mem[10][85] ), .IN4(n6776), .Q(n4066)
          );
   AO22X1 U3131 (.IN1(n7194), .IN2(n2505), .IN3(\key_mem[11][85] ), .IN4(n7189), .Q(n4067)
          );
   AO22X1 U3132 (.IN1(n6832), .IN2(n2505), .IN3(\key_mem[12][85] ), .IN4(n6839), .Q(n4068)
          );
   AO22X1 U3133 (.IN1(n7173), .IN2(n2505), .IN3(\key_mem[13][85] ), .IN4(n7168), .Q(n4069)
          );
   AO22X1 U3134 (.IN1(n7158), .IN2(n2505), .IN3(\key_mem[14][85] ), .IN4(n7149), .Q(n4070)
          );
   AO221X1 U3135 (.IN1(n7129), .IN2(n2506), .IN3(key[213]), .IN4(n7292), .IN5(n2507), .Q(
          n2505));
   AO222X1 U3136 (.IN1(n7115), .IN2(n2508), .IN3(key[85]), .IN4(n7074), .IN5(n7041), .IN6(
          n2509), .Q(n2507));
   AO22X1 U3137 (.IN1(n7298), .IN2(n2510), .IN3(\key_mem[0][84] ), .IN4(n6935), .Q(n4071)
          );
   AO22X1 U3138 (.IN1(n6813), .IN2(n2510), .IN3(\key_mem[1][84] ), .IN4(n6816), .Q(n4072)
          );
   AO22X1 U3139 (.IN1(n6857), .IN2(n2510), .IN3(\key_mem[2][84] ), .IN4(n6845), .Q(n4073)
          );
   AO22X1 U3140 (.IN1(n6873), .IN2(n2510), .IN3(\key_mem[3][84] ), .IN4(n6866), .Q(n4074)
          );
   AO22X1 U3141 (.IN1(n7286), .IN2(n2510), .IN3(\key_mem[4][84] ), .IN4(n6918), .Q(n4075)
          );
   AO22X1 U3142 (.IN1(n7275), .IN2(n2510), .IN3(\key_mem[5][84] ), .IN4(n7269), .Q(n4076)
          );
   AO22X1 U3143 (.IN1(n7017), .IN2(n2510), .IN3(\key_mem[6][84] ), .IN4(n7256), .Q(n4077)
          );
   AO22X1 U3144 (.IN1(n7013), .IN2(n2510), .IN3(\key_mem[7][84] ), .IN4(n7235), .Q(n4078)
          );
   AO22X1 U3145 (.IN1(n6757), .IN2(n2510), .IN3(\key_mem[8][84] ), .IN4(n6718), .Q(n4079)
          );
   AO22X1 U3146 (.IN1(n7219), .IN2(n2510), .IN3(\key_mem[9][84] ), .IN4(n7214), .Q(n4080)
          );
   AO22X1 U3147 (.IN1(n6804), .IN2(n2510), .IN3(\key_mem[10][84] ), .IN4(n6765), .Q(n4081)
          );
   AO22X1 U3148 (.IN1(n7195), .IN2(n2510), .IN3(\key_mem[11][84] ), .IN4(n7190), .Q(n4082)
          );
   AO22X1 U3149 (.IN1(n6829), .IN2(n2510), .IN3(\key_mem[12][84] ), .IN4(n6983), .Q(n4083)
          );
   AO22X1 U3150 (.IN1(n7174), .IN2(n2510), .IN3(\key_mem[13][84] ), .IN4(n7169), .Q(n4084)
          );
   AO22X1 U3151 (.IN1(n7159), .IN2(n2510), .IN3(\key_mem[14][84] ), .IN4(n7156), .Q(n4085)
          );
   AO221X1 U3152 (.IN1(n7129), .IN2(n2511), .IN3(key[212]), .IN4(n7294), .IN5(n2512), .Q(
          n2510));
   AO222X1 U3153 (.IN1(n7115), .IN2(n2513), .IN3(key[84]), .IN4(n7074), .IN5(n7041), .IN6(
          n2514), .Q(n2512));
   AO22X1 U3154 (.IN1(n7297), .IN2(n2515), .IN3(\key_mem[0][83] ), .IN4(n6934), .Q(n4086)
          );
   AO22X1 U3155 (.IN1(n6813), .IN2(n2515), .IN3(\key_mem[1][83] ), .IN4(n6818), .Q(n4087)
          );
   AO22X1 U3156 (.IN1(n6854), .IN2(n2515), .IN3(\key_mem[2][83] ), .IN4(n6843), .Q(n4088)
          );
   AO22X1 U3157 (.IN1(n6874), .IN2(n2515), .IN3(\key_mem[3][83] ), .IN4(n6865), .Q(n4089)
          );
   AO22X1 U3158 (.IN1(n6886), .IN2(n2515), .IN3(\key_mem[4][83] ), .IN4(n6923), .Q(n4090)
          );
   AO22X1 U3159 (.IN1(n7275), .IN2(n2515), .IN3(\key_mem[5][83] ), .IN4(n7272), .Q(n4091)
          );
   AO22X1 U3160 (.IN1(n7016), .IN2(n2515), .IN3(\key_mem[6][83] ), .IN4(n7255), .Q(n4092)
          );
   AO22X1 U3161 (.IN1(n7247), .IN2(n2515), .IN3(\key_mem[7][83] ), .IN4(n7236), .Q(n4093)
          );
   AO22X1 U3162 (.IN1(n6758), .IN2(n2515), .IN3(\key_mem[8][83] ), .IN4(n6724), .Q(n4094)
          );
   AO22X1 U3163 (.IN1(n7219), .IN2(n2515), .IN3(\key_mem[9][83] ), .IN4(n7216), .Q(n4095)
          );
   AO22X1 U3164 (.IN1(n6805), .IN2(n2515), .IN3(\key_mem[10][83] ), .IN4(n6771), .Q(n4096)
          );
   AO22X1 U3165 (.IN1(n7195), .IN2(n2515), .IN3(\key_mem[11][83] ), .IN4(n7192), .Q(n4097)
          );
   AO22X1 U3166 (.IN1(n6829), .IN2(n2515), .IN3(\key_mem[12][83] ), .IN4(n2289), .Q(n4098)
          );
   AO22X1 U3167 (.IN1(n7174), .IN2(n2515), .IN3(\key_mem[13][83] ), .IN4(n7171), .Q(n4099)
          );
   AO22X1 U3168 (.IN1(n6972), .IN2(n2515), .IN3(\key_mem[14][83] ), .IN4(n7165), .Q(n4100)
          );
   AO221X1 U3169 (.IN1(n7129), .IN2(n2516), .IN3(key[211]), .IN4(n7292), .IN5(n2517), .Q(
          n2515));
   AO222X1 U3170 (.IN1(n7115), .IN2(n2518), .IN3(key[83]), .IN4(n7074), .IN5(n7041), .IN6(
          n2519), .Q(n2517));
   AO22X1 U3171 (.IN1(n7296), .IN2(n2520), .IN3(\key_mem[0][82] ), .IN4(n6934), .Q(n4101)
          );
   AO22X1 U3172 (.IN1(n6809), .IN2(n2520), .IN3(\key_mem[1][82] ), .IN4(n6819), .Q(n4102)
          );
   AO22X1 U3173 (.IN1(n6855), .IN2(n2520), .IN3(\key_mem[2][82] ), .IN4(n6848), .Q(n4103)
          );
   AO22X1 U3174 (.IN1(n6873), .IN2(n2520), .IN3(\key_mem[3][82] ), .IN4(n6868), .Q(n4104)
          );
   AO22X1 U3175 (.IN1(n6889), .IN2(n2520), .IN3(\key_mem[4][82] ), .IN4(n6915), .Q(n4105)
          );
   AO22X1 U3176 (.IN1(n7019), .IN2(n2520), .IN3(\key_mem[5][82] ), .IN4(n7267), .Q(n4106)
          );
   AO22X1 U3177 (.IN1(n7260), .IN2(n2520), .IN3(\key_mem[6][82] ), .IN4(n7252), .Q(n4107)
          );
   AO22X1 U3178 (.IN1(n7247), .IN2(n2520), .IN3(\key_mem[7][82] ), .IN4(n7237), .Q(n4108)
          );
   AO22X1 U3179 (.IN1(n6755), .IN2(n2520), .IN3(\key_mem[8][82] ), .IN4(n6721), .Q(n4109)
          );
   AO22X1 U3180 (.IN1(n7008), .IN2(n2520), .IN3(\key_mem[9][82] ), .IN4(n7211), .Q(n4110)
          );
   AO22X1 U3181 (.IN1(n6802), .IN2(n2520), .IN3(\key_mem[10][82] ), .IN4(n6768), .Q(n4111)
          );
   AO22X1 U3182 (.IN1(n7003), .IN2(n2520), .IN3(\key_mem[11][82] ), .IN4(n7187), .Q(n4112)
          );
   AO22X1 U3183 (.IN1(n7001), .IN2(n2520), .IN3(\key_mem[12][82] ), .IN4(n7185), .Q(n4113)
          );
   AO22X1 U3184 (.IN1(n6998), .IN2(n2520), .IN3(\key_mem[13][82] ), .IN4(n7166), .Q(n4114)
          );
   AO22X1 U3185 (.IN1(n7163), .IN2(n2520), .IN3(\key_mem[14][82] ), .IN4(n6994), .Q(n4115)
          );
   AO221X1 U3186 (.IN1(n7129), .IN2(n2521), .IN3(key[210]), .IN4(n7291), .IN5(n2522), .Q(
          n2520));
   AO222X1 U3187 (.IN1(n7114), .IN2(n2523), .IN3(key[82]), .IN4(n7074), .IN5(n7041), .IN6(
          n2524), .Q(n2522));
   AO22X1 U3188 (.IN1(n7295), .IN2(n2525), .IN3(\key_mem[0][81] ), .IN4(n6934), .Q(n4116)
          );
   AO22X1 U3189 (.IN1(n6811), .IN2(n2525), .IN3(\key_mem[1][81] ), .IN4(n6817), .Q(n4117)
          );
   AO22X1 U3190 (.IN1(n6857), .IN2(n2525), .IN3(\key_mem[2][81] ), .IN4(n6850), .Q(n4118)
          );
   AO22X1 U3191 (.IN1(n6807), .IN2(n2525), .IN3(\key_mem[3][81] ), .IN4(n6860), .Q(n4119)
          );
   AO22X1 U3192 (.IN1(n6922), .IN2(n2525), .IN3(\key_mem[4][81] ), .IN4(n6923), .Q(n4120)
          );
   AO22X1 U3193 (.IN1(n7283), .IN2(n2525), .IN3(\key_mem[5][81] ), .IN4(n7273), .Q(n4121)
          );
   AO22X1 U3194 (.IN1(n7016), .IN2(n2525), .IN3(\key_mem[6][81] ), .IN4(n7253), .Q(n4122)
          );
   AO22X1 U3195 (.IN1(n7249), .IN2(n2525), .IN3(\key_mem[7][81] ), .IN4(n7238), .Q(n4123)
          );
   AO22X1 U3196 (.IN1(n6756), .IN2(n2525), .IN3(\key_mem[8][81] ), .IN4(n6717), .Q(n4124)
          );
   AO22X1 U3197 (.IN1(n7227), .IN2(n2525), .IN3(\key_mem[9][81] ), .IN4(n7217), .Q(n4125)
          );
   AO22X1 U3198 (.IN1(n6803), .IN2(n2525), .IN3(\key_mem[10][81] ), .IN4(n6764), .Q(n4126)
          );
   AO22X1 U3199 (.IN1(n7203), .IN2(n2525), .IN3(\key_mem[11][81] ), .IN4(n7193), .Q(n4127)
          );
   AO22X1 U3200 (.IN1(n6827), .IN2(n2525), .IN3(\key_mem[12][81] ), .IN4(n6982), .Q(n4128)
          );
   AO22X1 U3201 (.IN1(n7182), .IN2(n2525), .IN3(\key_mem[13][81] ), .IN4(n7172), .Q(n4129)
          );
   AO22X1 U3202 (.IN1(n7162), .IN2(n2525), .IN3(\key_mem[14][81] ), .IN4(n7151), .Q(n4130)
          );
   AO221X1 U3203 (.IN1(n7129), .IN2(n2526), .IN3(key[209]), .IN4(n7299), .IN5(n2527), .Q(
          n2525));
   AO222X1 U3204 (.IN1(n7114), .IN2(n2528), .IN3(key[81]), .IN4(n7074), .IN5(n7041), .IN6(
          n2529), .Q(n2527));
   AO22X1 U3205 (.IN1(n7304), .IN2(n2530), .IN3(\key_mem[0][80] ), .IN4(n6934), .Q(n4131)
          );
   AO22X1 U3206 (.IN1(n6926), .IN2(n2530), .IN3(\key_mem[1][80] ), .IN4(n6818), .Q(n4132)
          );
   AO22X1 U3207 (.IN1(n6853), .IN2(n2530), .IN3(\key_mem[2][80] ), .IN4(n6849), .Q(n4133)
          );
   AO22X1 U3208 (.IN1(n6989), .IN2(n2530), .IN3(\key_mem[3][80] ), .IN4(n6862), .Q(n4134)
          );
   AO22X1 U3209 (.IN1(n6922), .IN2(n2530), .IN3(\key_mem[4][80] ), .IN4(n7021), .Q(n4135)
          );
   AO22X1 U3210 (.IN1(n6973), .IN2(n2530), .IN3(\key_mem[5][80] ), .IN4(n7271), .Q(n4136)
          );
   AO22X1 U3211 (.IN1(n7016), .IN2(n2530), .IN3(\key_mem[6][80] ), .IN4(n7259), .Q(n4137)
          );
   AO22X1 U3212 (.IN1(n7248), .IN2(n2530), .IN3(\key_mem[7][80] ), .IN4(n7239), .Q(n4138)
          );
   AO22X1 U3213 (.IN1(n6757), .IN2(n2530), .IN3(\key_mem[8][80] ), .IN4(n6743), .Q(n4139)
          );
   AO22X1 U3214 (.IN1(n7218), .IN2(n2530), .IN3(\key_mem[9][80] ), .IN4(n7215), .Q(n4140)
          );
   AO22X1 U3215 (.IN1(n6804), .IN2(n2530), .IN3(\key_mem[10][80] ), .IN4(n6790), .Q(n4141)
          );
   AO22X1 U3216 (.IN1(n7194), .IN2(n2530), .IN3(\key_mem[11][80] ), .IN4(n7191), .Q(n4142)
          );
   AO22X1 U3217 (.IN1(n7183), .IN2(n2530), .IN3(\key_mem[12][80] ), .IN4(n6985), .Q(n4143)
          );
   AO22X1 U3218 (.IN1(n7173), .IN2(n2530), .IN3(\key_mem[13][80] ), .IN4(n7170), .Q(n4144)
          );
   AO22X1 U3219 (.IN1(n7163), .IN2(n2530), .IN3(\key_mem[14][80] ), .IN4(n7152), .Q(n4145)
          );
   AO221X1 U3220 (.IN1(n7129), .IN2(n2531), .IN3(key[208]), .IN4(n7298), .IN5(n2532), .Q(
          n2530));
   AO222X1 U3221 (.IN1(n7114), .IN2(n2533), .IN3(key[80]), .IN4(n7074), .IN5(n7041), .IN6(
          n2534), .Q(n2532));
   AO22X1 U3222 (.IN1(n7303), .IN2(n2535), .IN3(\key_mem[0][79] ), .IN4(n6934), .Q(n4146)
          );
   AO22X1 U3223 (.IN1(n6808), .IN2(n2535), .IN3(\key_mem[1][79] ), .IN4(n6822), .Q(n4147)
          );
   AO22X1 U3224 (.IN1(n6858), .IN2(n2535), .IN3(\key_mem[2][79] ), .IN4(n6847), .Q(n4148)
          );
   AO22X1 U3225 (.IN1(n6807), .IN2(n2535), .IN3(\key_mem[3][79] ), .IN4(n6863), .Q(n4149)
          );
   AO22X1 U3226 (.IN1(n6924), .IN2(n2535), .IN3(\key_mem[4][79] ), .IN4(n7284), .Q(n4150)
          );
   AO22X1 U3227 (.IN1(n7274), .IN2(n2535), .IN3(\key_mem[5][79] ), .IN4(n7272), .Q(n4151)
          );
   AO22X1 U3228 (.IN1(n7016), .IN2(n2535), .IN3(\key_mem[6][79] ), .IN4(n7251), .Q(n4152)
          );
   AO22X1 U3229 (.IN1(n7247), .IN2(n2535), .IN3(\key_mem[7][79] ), .IN4(n7240), .Q(n4153)
          );
   AO22X1 U3230 (.IN1(n6758), .IN2(n2535), .IN3(\key_mem[8][79] ), .IN4(n6745), .Q(n4154)
          );
   AO22X1 U3231 (.IN1(n6976), .IN2(n2535), .IN3(\key_mem[9][79] ), .IN4(n7216), .Q(n4155)
          );
   AO22X1 U3232 (.IN1(n6805), .IN2(n2535), .IN3(\key_mem[10][79] ), .IN4(n6792), .Q(n4156)
          );
   AO22X1 U3233 (.IN1(n6978), .IN2(n2535), .IN3(\key_mem[11][79] ), .IN4(n7192), .Q(n4157)
          );
   AO22X1 U3234 (.IN1(n6829), .IN2(n2535), .IN3(\key_mem[12][79] ), .IN4(n6830), .Q(n4158)
          );
   AO22X1 U3235 (.IN1(n6980), .IN2(n2535), .IN3(\key_mem[13][79] ), .IN4(n7171), .Q(n4159)
          );
   AO22X1 U3236 (.IN1(n7161), .IN2(n2535), .IN3(\key_mem[14][79] ), .IN4(n7153), .Q(n4160)
          );
   AO221X1 U3237 (.IN1(n7130), .IN2(n2536), .IN3(key[207]), .IN4(n7297), .IN5(n2537), .Q(
          n2535));
   AO222X1 U3238 (.IN1(n7114), .IN2(n2538), .IN3(key[79]), .IN4(n7075), .IN5(n7042), .IN6(
          n2539), .Q(n2537));
   AO22X1 U3239 (.IN1(n7302), .IN2(n2540), .IN3(\key_mem[0][78] ), .IN4(n6934), .Q(n4161)
          );
   AO22X1 U3240 (.IN1(n6926), .IN2(n2540), .IN3(\key_mem[1][78] ), .IN4(n6816), .Q(n4162)
          );
   AO22X1 U3241 (.IN1(n6854), .IN2(n2540), .IN3(\key_mem[2][78] ), .IN4(n6846), .Q(n4163)
          );
   AO22X1 U3242 (.IN1(n6989), .IN2(n2540), .IN3(\key_mem[3][78] ), .IN4(n6862), .Q(n4164)
          );
   AO22X1 U3243 (.IN1(n6889), .IN2(n2540), .IN3(\key_mem[4][78] ), .IN4(n6923), .Q(n4165)
          );
   AO22X1 U3244 (.IN1(n7275), .IN2(n2540), .IN3(\key_mem[5][78] ), .IN4(n7267), .Q(n4166)
          );
   AO22X1 U3245 (.IN1(n7262), .IN2(n2540), .IN3(\key_mem[6][78] ), .IN4(n7256), .Q(n4167)
          );
   AO22X1 U3246 (.IN1(n7246), .IN2(n2540), .IN3(\key_mem[7][78] ), .IN4(n7241), .Q(n4168)
          );
   AO22X1 U3247 (.IN1(n6748), .IN2(n2540), .IN3(\key_mem[8][78] ), .IN4(n6746), .Q(n4169)
          );
   AO22X1 U3248 (.IN1(n7223), .IN2(n2540), .IN3(\key_mem[9][78] ), .IN4(n7217), .Q(n4170)
          );
   AO22X1 U3249 (.IN1(n6795), .IN2(n2540), .IN3(\key_mem[10][78] ), .IN4(n6793), .Q(n4171)
          );
   AO22X1 U3250 (.IN1(n7199), .IN2(n2540), .IN3(\key_mem[11][78] ), .IN4(n7193), .Q(n4172)
          );
   AO22X1 U3251 (.IN1(n6832), .IN2(n2540), .IN3(\key_mem[12][78] ), .IN4(n6982), .Q(n4173)
          );
   AO22X1 U3252 (.IN1(n7178), .IN2(n2540), .IN3(\key_mem[13][78] ), .IN4(n7172), .Q(n4174)
          );
   AO22X1 U3253 (.IN1(n7160), .IN2(n2540), .IN3(\key_mem[14][78] ), .IN4(n7154), .Q(n4175)
          );
   AO221X1 U3254 (.IN1(n7130), .IN2(n2541), .IN3(key[206]), .IN4(n7293), .IN5(n2542), .Q(
          n2540));
   AO222X1 U3255 (.IN1(n7114), .IN2(n2543), .IN3(key[78]), .IN4(n7075), .IN5(n7042), .IN6(
          n2544), .Q(n2542));
   AO22X1 U3256 (.IN1(n7301), .IN2(n2545), .IN3(\key_mem[0][77] ), .IN4(n6934), .Q(n4176)
          );
   AO22X1 U3257 (.IN1(n6812), .IN2(n2545), .IN3(\key_mem[1][77] ), .IN4(n6823), .Q(n4177)
          );
   AO22X1 U3258 (.IN1(n6854), .IN2(n2545), .IN3(\key_mem[2][77] ), .IN4(n6859), .Q(n4178)
          );
   AO22X1 U3259 (.IN1(n6872), .IN2(n2545), .IN3(\key_mem[3][77] ), .IN4(n6868), .Q(n4179)
          );
   AO22X1 U3260 (.IN1(n6886), .IN2(n2545), .IN3(\key_mem[4][77] ), .IN4(n7285), .Q(n4180)
          );
   AO22X1 U3261 (.IN1(n6974), .IN2(n2545), .IN3(\key_mem[5][77] ), .IN4(n7282), .Q(n4181)
          );
   AO22X1 U3262 (.IN1(n7263), .IN2(n2545), .IN3(\key_mem[6][77] ), .IN4(n7254), .Q(n4182)
          );
   AO22X1 U3263 (.IN1(n7245), .IN2(n2545), .IN3(\key_mem[7][77] ), .IN4(n7235), .Q(n4183)
          );
   AO22X1 U3264 (.IN1(n6748), .IN2(n2545), .IN3(\key_mem[8][77] ), .IN4(n6731), .Q(n4184)
          );
   AO22X1 U3265 (.IN1(n6975), .IN2(n2545), .IN3(\key_mem[9][77] ), .IN4(n7226), .Q(n4185)
          );
   AO22X1 U3266 (.IN1(n6795), .IN2(n2545), .IN3(\key_mem[10][77] ), .IN4(n6778), .Q(n4186)
          );
   AO22X1 U3267 (.IN1(n6977), .IN2(n2545), .IN3(\key_mem[11][77] ), .IN4(n7202), .Q(n4187)
          );
   AO22X1 U3268 (.IN1(n6831), .IN2(n2545), .IN3(\key_mem[12][77] ), .IN4(n6833), .Q(n4188)
          );
   AO22X1 U3269 (.IN1(n6979), .IN2(n2545), .IN3(\key_mem[13][77] ), .IN4(n7181), .Q(n4189)
          );
   AO22X1 U3270 (.IN1(n7161), .IN2(n2545), .IN3(\key_mem[14][77] ), .IN4(n7155), .Q(n4190)
          );
   AO221X1 U3271 (.IN1(n7130), .IN2(n2546), .IN3(key[205]), .IN4(n7291), .IN5(n2547), .Q(
          n2545));
   AO222X1 U3272 (.IN1(n7114), .IN2(n2548), .IN3(key[77]), .IN4(n7075), .IN5(n7042), .IN6(
          n2549), .Q(n2547));
   AO22X1 U3273 (.IN1(n7311), .IN2(n2550), .IN3(\key_mem[0][76] ), .IN4(n6934), .Q(n4191)
          );
   AO22X1 U3274 (.IN1(n6808), .IN2(n2550), .IN3(\key_mem[1][76] ), .IN4(n6821), .Q(n4192)
          );
   AO22X1 U3275 (.IN1(n6856), .IN2(n2550), .IN3(\key_mem[2][76] ), .IN4(n6842), .Q(n4193)
          );
   AO22X1 U3276 (.IN1(n6869), .IN2(n2550), .IN3(\key_mem[3][76] ), .IN4(n6867), .Q(n4194)
          );
   AO22X1 U3277 (.IN1(n6887), .IN2(n2550), .IN3(\key_mem[4][76] ), .IN4(n6925), .Q(n4195)
          );
   AO22X1 U3278 (.IN1(n7279), .IN2(n2550), .IN3(\key_mem[5][76] ), .IN4(n7273), .Q(n4196)
          );
   AO22X1 U3279 (.IN1(n7261), .IN2(n2550), .IN3(\key_mem[6][76] ), .IN4(n7258), .Q(n4197)
          );
   AO22X1 U3280 (.IN1(n7244), .IN2(n2550), .IN3(\key_mem[7][76] ), .IN4(n7235), .Q(n4198)
          );
   AO22X1 U3281 (.IN1(n6749), .IN2(n2550), .IN3(\key_mem[8][76] ), .IN4(n6733), .Q(n4199)
          );
   AO22X1 U3282 (.IN1(n7219), .IN2(n2550), .IN3(\key_mem[9][76] ), .IN4(n7217), .Q(n4200)
          );
   AO22X1 U3283 (.IN1(n6796), .IN2(n2550), .IN3(\key_mem[10][76] ), .IN4(n6780), .Q(n4201)
          );
   AO22X1 U3284 (.IN1(n7195), .IN2(n2550), .IN3(\key_mem[11][76] ), .IN4(n7193), .Q(n4202)
          );
   AO22X1 U3285 (.IN1(n6826), .IN2(n2550), .IN3(\key_mem[12][76] ), .IN4(n6981), .Q(n4203)
          );
   AO22X1 U3286 (.IN1(n7174), .IN2(n2550), .IN3(\key_mem[13][76] ), .IN4(n7172), .Q(n4204)
          );
   AO22X1 U3287 (.IN1(n6996), .IN2(n2550), .IN3(\key_mem[14][76] ), .IN4(n7147), .Q(n4205)
          );
   AO221X1 U3288 (.IN1(n7130), .IN2(n2551), .IN3(key[204]), .IN4(n7290), .IN5(n2552), .Q(
          n2550));
   AO222X1 U3289 (.IN1(n7114), .IN2(n2553), .IN3(key[76]), .IN4(n7075), .IN5(n7042), .IN6(
          n2554), .Q(n2552));
   AO22X1 U3290 (.IN1(n7300), .IN2(n2555), .IN3(\key_mem[0][75] ), .IN4(n6934), .Q(n4206)
          );
   AO22X1 U3291 (.IN1(n6926), .IN2(n2555), .IN3(\key_mem[1][75] ), .IN4(n6815), .Q(n4207)
          );
   AO22X1 U3292 (.IN1(n6988), .IN2(n2555), .IN3(\key_mem[2][75] ), .IN4(n6847), .Q(n4208)
          );
   AO22X1 U3293 (.IN1(n6870), .IN2(n2555), .IN3(\key_mem[3][75] ), .IN4(n6876), .Q(n4209)
          );
   AO22X1 U3294 (.IN1(n6922), .IN2(n2555), .IN3(\key_mem[4][75] ), .IN4(n6915), .Q(n4210)
          );
   AO22X1 U3295 (.IN1(n7277), .IN2(n2555), .IN3(\key_mem[5][75] ), .IN4(n2282), .Q(n4211)
          );
   AO22X1 U3296 (.IN1(n6969), .IN2(n2555), .IN3(\key_mem[6][75] ), .IN4(n7256), .Q(n4212)
          );
   AO22X1 U3297 (.IN1(n7249), .IN2(n2555), .IN3(\key_mem[7][75] ), .IN4(n7241), .Q(n4213)
          );
   AO22X1 U3298 (.IN1(n6750), .IN2(n2555), .IN3(\key_mem[8][75] ), .IN4(n6734), .Q(n4214)
          );
   AO22X1 U3299 (.IN1(n7221), .IN2(n2555), .IN3(\key_mem[9][75] ), .IN4(n2286), .Q(n4215)
          );
   AO22X1 U3300 (.IN1(n6797), .IN2(n2555), .IN3(\key_mem[10][75] ), .IN4(n6781), .Q(n4216)
          );
   AO22X1 U3301 (.IN1(n7197), .IN2(n2555), .IN3(\key_mem[11][75] ), .IN4(n2288), .Q(n4217)
          );
   AO22X1 U3302 (.IN1(n6826), .IN2(n2555), .IN3(\key_mem[12][75] ), .IN4(n7000), .Q(n4218)
          );
   AO22X1 U3303 (.IN1(n7176), .IN2(n2555), .IN3(\key_mem[13][75] ), .IN4(n2290), .Q(n4219)
          );
   AO22X1 U3304 (.IN1(n7162), .IN2(n2555), .IN3(\key_mem[14][75] ), .IN4(n7165), .Q(n4220)
          );
   AO221X1 U3305 (.IN1(n7130), .IN2(n2556), .IN3(key[203]), .IN4(n7298), .IN5(n2557), .Q(
          n2555));
   AO222X1 U3306 (.IN1(n7114), .IN2(n2558), .IN3(key[75]), .IN4(n7075), .IN5(n7042), .IN6(
          n2559), .Q(n2557));
   AO22X1 U3307 (.IN1(n7292), .IN2(n2560), .IN3(\key_mem[0][74] ), .IN4(n6934), .Q(n4221)
          );
   AO22X1 U3308 (.IN1(n6926), .IN2(n2560), .IN3(\key_mem[1][74] ), .IN4(n6817), .Q(n4222)
          );
   AO22X1 U3309 (.IN1(n6852), .IN2(n2560), .IN3(\key_mem[2][74] ), .IN4(n6859), .Q(n4223)
          );
   AO22X1 U3310 (.IN1(n6806), .IN2(n2560), .IN3(\key_mem[3][74] ), .IN4(n6877), .Q(n4224)
          );
   AO22X1 U3311 (.IN1(n6922), .IN2(n2560), .IN3(\key_mem[4][74] ), .IN4(n7284), .Q(n4225)
          );
   AO22X1 U3312 (.IN1(n7276), .IN2(n2560), .IN3(\key_mem[5][74] ), .IN4(n7281), .Q(n4226)
          );
   AO22X1 U3313 (.IN1(n6970), .IN2(n2560), .IN3(\key_mem[6][74] ), .IN4(n7254), .Q(n4227)
          );
   AO22X1 U3314 (.IN1(n7246), .IN2(n2560), .IN3(\key_mem[7][74] ), .IN4(n7239), .Q(n4228)
          );
   AO22X1 U3315 (.IN1(n6748), .IN2(n2560), .IN3(\key_mem[8][74] ), .IN4(n6721), .Q(n4229)
          );
   AO22X1 U3316 (.IN1(n7220), .IN2(n2560), .IN3(\key_mem[9][74] ), .IN4(n7225), .Q(n4230)
          );
   AO22X1 U3317 (.IN1(n6795), .IN2(n2560), .IN3(\key_mem[10][74] ), .IN4(n6768), .Q(n4231)
          );
   AO22X1 U3318 (.IN1(n7196), .IN2(n2560), .IN3(\key_mem[11][74] ), .IN4(n7201), .Q(n4232)
          );
   AO22X1 U3319 (.IN1(n6837), .IN2(n2560), .IN3(\key_mem[12][74] ), .IN4(n6834), .Q(n4233)
          );
   AO22X1 U3320 (.IN1(n7175), .IN2(n2560), .IN3(\key_mem[13][74] ), .IN4(n7180), .Q(n4234)
          );
   AO22X1 U3321 (.IN1(n6996), .IN2(n2560), .IN3(\key_mem[14][74] ), .IN4(n7153), .Q(n4235)
          );
   AO221X1 U3322 (.IN1(n7130), .IN2(n2561), .IN3(key[202]), .IN4(n7297), .IN5(n2562), .Q(
          n2560));
   AO222X1 U3323 (.IN1(n7114), .IN2(n2563), .IN3(key[74]), .IN4(n7075), .IN5(n7042), .IN6(
          n2564), .Q(n2562));
   AO22X1 U3324 (.IN1(n7295), .IN2(n2565), .IN3(\key_mem[0][73] ), .IN4(n6934), .Q(n4236)
          );
   AO22X1 U3325 (.IN1(n6809), .IN2(n2565), .IN3(\key_mem[1][73] ), .IN4(n6818), .Q(n4237)
          );
   AO22X1 U3326 (.IN1(n6854), .IN2(n2565), .IN3(\key_mem[2][73] ), .IN4(n6844), .Q(n4238)
          );
   AO22X1 U3327 (.IN1(n6871), .IN2(n2565), .IN3(\key_mem[3][73] ), .IN4(n6863), .Q(n4239)
          );
   AO22X1 U3328 (.IN1(n6990), .IN2(n2565), .IN3(\key_mem[4][73] ), .IN4(n6925), .Q(n4240)
          );
   AO22X1 U3329 (.IN1(n7277), .IN2(n2565), .IN3(\key_mem[5][73] ), .IN4(n7273), .Q(n4241)
          );
   AO22X1 U3330 (.IN1(n7265), .IN2(n2565), .IN3(\key_mem[6][73] ), .IN4(n2283), .Q(n4242)
          );
   AO22X1 U3331 (.IN1(n7246), .IN2(n2565), .IN3(\key_mem[7][73] ), .IN4(n7242), .Q(n4243)
          );
   AO22X1 U3332 (.IN1(n6749), .IN2(n2565), .IN3(\key_mem[8][73] ), .IN4(n6722), .Q(n4244)
          );
   AO22X1 U3333 (.IN1(n7221), .IN2(n2565), .IN3(\key_mem[9][73] ), .IN4(n7217), .Q(n4245)
          );
   AO22X1 U3334 (.IN1(n6796), .IN2(n2565), .IN3(\key_mem[10][73] ), .IN4(n6769), .Q(n4246)
          );
   AO22X1 U3335 (.IN1(n7197), .IN2(n2565), .IN3(\key_mem[11][73] ), .IN4(n7193), .Q(n4247)
          );
   AO22X1 U3336 (.IN1(n6827), .IN2(n2565), .IN3(\key_mem[12][73] ), .IN4(n7184), .Q(n4248)
          );
   AO22X1 U3337 (.IN1(n7176), .IN2(n2565), .IN3(\key_mem[13][73] ), .IN4(n7172), .Q(n4249)
          );
   AO22X1 U3338 (.IN1(n6995), .IN2(n2565), .IN3(\key_mem[14][73] ), .IN4(n7154), .Q(n4250)
          );
   AO221X1 U3339 (.IN1(n7130), .IN2(n2566), .IN3(key[201]), .IN4(n7295), .IN5(n2567), .Q(
          n2565));
   AO222X1 U3340 (.IN1(n7114), .IN2(n2568), .IN3(key[73]), .IN4(n7075), .IN5(n7042), .IN6(
          n2569), .Q(n2567));
   AO22X1 U3341 (.IN1(n7304), .IN2(n2570), .IN3(\key_mem[0][72] ), .IN4(n6934), .Q(n4251)
          );
   AO22X1 U3342 (.IN1(n6810), .IN2(n2570), .IN3(\key_mem[1][72] ), .IN4(n6817), .Q(n4252)
          );
   AO22X1 U3343 (.IN1(n6857), .IN2(n2570), .IN3(\key_mem[2][72] ), .IN4(n6845), .Q(n4253)
          );
   AO22X1 U3344 (.IN1(n6806), .IN2(n2570), .IN3(\key_mem[3][72] ), .IN4(n6876), .Q(n4254)
          );
   AO22X1 U3345 (.IN1(n7286), .IN2(n2570), .IN3(\key_mem[4][72] ), .IN4(n6923), .Q(n4255)
          );
   AO22X1 U3346 (.IN1(n7276), .IN2(n2570), .IN3(\key_mem[5][72] ), .IN4(n7273), .Q(n4256)
          );
   AO22X1 U3347 (.IN1(n7260), .IN2(n2570), .IN3(\key_mem[6][72] ), .IN4(n7015), .Q(n4257)
          );
   AO22X1 U3348 (.IN1(n7250), .IN2(n2570), .IN3(\key_mem[7][72] ), .IN4(n7238), .Q(n4258)
          );
   AO22X1 U3349 (.IN1(n6749), .IN2(n2570), .IN3(\key_mem[8][72] ), .IN4(n6717), .Q(n4259)
          );
   AO22X1 U3350 (.IN1(n7220), .IN2(n2570), .IN3(\key_mem[9][72] ), .IN4(n7217), .Q(n4260)
          );
   AO22X1 U3351 (.IN1(n6796), .IN2(n2570), .IN3(\key_mem[10][72] ), .IN4(n6764), .Q(n4261)
          );
   AO22X1 U3352 (.IN1(n7196), .IN2(n2570), .IN3(\key_mem[11][72] ), .IN4(n7193), .Q(n4262)
          );
   AO22X1 U3353 (.IN1(n7186), .IN2(n2570), .IN3(\key_mem[12][72] ), .IN4(n6830), .Q(n4263)
          );
   AO22X1 U3354 (.IN1(n7175), .IN2(n2570), .IN3(\key_mem[13][72] ), .IN4(n7172), .Q(n4264)
          );
   AO22X1 U3355 (.IN1(n6992), .IN2(n2570), .IN3(\key_mem[14][72] ), .IN4(n6994), .Q(n4265)
          );
   AO221X1 U3356 (.IN1(n7130), .IN2(n2571), .IN3(key[200]), .IN4(n7304), .IN5(n2572), .Q(
          n2570));
   AO222X1 U3357 (.IN1(n7114), .IN2(n2573), .IN3(key[72]), .IN4(n7075), .IN5(n7042), .IN6(
          n2574), .Q(n2572));
   AO22X1 U3358 (.IN1(n7303), .IN2(n2575), .IN3(\key_mem[0][71] ), .IN4(n6933), .Q(n4266)
          );
   AO22X1 U3359 (.IN1(n6808), .IN2(n2575), .IN3(\key_mem[1][71] ), .IN4(n6814), .Q(n4267)
          );
   AO22X1 U3360 (.IN1(n6852), .IN2(n2575), .IN3(\key_mem[2][71] ), .IN4(n6847), .Q(n4268)
          );
   AO22X1 U3361 (.IN1(n6869), .IN2(n2575), .IN3(\key_mem[3][71] ), .IN4(n6862), .Q(n4269)
          );
   AO22X1 U3362 (.IN1(n6887), .IN2(n2575), .IN3(\key_mem[4][71] ), .IN4(n7284), .Q(n4270)
          );
   AO22X1 U3363 (.IN1(n7276), .IN2(n2575), .IN3(\key_mem[5][71] ), .IN4(n7268), .Q(n4271)
          );
   AO22X1 U3364 (.IN1(n7261), .IN2(n2575), .IN3(\key_mem[6][71] ), .IN4(n7251), .Q(n4272)
          );
   AO22X1 U3365 (.IN1(n7014), .IN2(n2575), .IN3(\key_mem[7][71] ), .IN4(n7012), .Q(n4273)
          );
   AO22X1 U3366 (.IN1(n6756), .IN2(n2575), .IN3(\key_mem[8][71] ), .IN4(n6724), .Q(n4274)
          );
   AO22X1 U3367 (.IN1(n7220), .IN2(n2575), .IN3(\key_mem[9][71] ), .IN4(n7216), .Q(n4275)
          );
   AO22X1 U3368 (.IN1(n6803), .IN2(n2575), .IN3(\key_mem[10][71] ), .IN4(n6771), .Q(n4276)
          );
   AO22X1 U3369 (.IN1(n7196), .IN2(n2575), .IN3(\key_mem[11][71] ), .IN4(n7192), .Q(n4277)
          );
   AO22X1 U3370 (.IN1(n6986), .IN2(n2575), .IN3(\key_mem[12][71] ), .IN4(n6836), .Q(n4278)
          );
   AO22X1 U3371 (.IN1(n7175), .IN2(n2575), .IN3(\key_mem[13][71] ), .IN4(n7171), .Q(n4279)
          );
   AO22X1 U3372 (.IN1(n7160), .IN2(n2575), .IN3(\key_mem[14][71] ), .IN4(n7157), .Q(n4280)
          );
   AO221X1 U3373 (.IN1(n7130), .IN2(n2576), .IN3(key[199]), .IN4(n7302), .IN5(n2577), .Q(
          n2575));
   AO222X1 U3374 (.IN1(n7114), .IN2(n2578), .IN3(key[71]), .IN4(n7075), .IN5(n7042), .IN6(
          n2579), .Q(n2577));
   AO22X1 U3375 (.IN1(n7302), .IN2(n2580), .IN3(\key_mem[0][70] ), .IN4(n6933), .Q(n4281)
          );
   AO22X1 U3376 (.IN1(n6809), .IN2(n2580), .IN3(\key_mem[1][70] ), .IN4(n6818), .Q(n4282)
          );
   AO22X1 U3377 (.IN1(n6852), .IN2(n2580), .IN3(\key_mem[2][70] ), .IN4(n6842), .Q(n4283)
          );
   AO22X1 U3378 (.IN1(n6869), .IN2(n2580), .IN3(\key_mem[3][70] ), .IN4(n6866), .Q(n4284)
          );
   AO22X1 U3379 (.IN1(n7022), .IN2(n2580), .IN3(\key_mem[4][70] ), .IN4(n6918), .Q(n4285)
          );
   AO22X1 U3380 (.IN1(n7279), .IN2(n2580), .IN3(\key_mem[5][70] ), .IN4(n7268), .Q(n4286)
          );
   AO22X1 U3381 (.IN1(n7260), .IN2(n2580), .IN3(\key_mem[6][70] ), .IN4(n7251), .Q(n4287)
          );
   AO22X1 U3382 (.IN1(n7247), .IN2(n2580), .IN3(\key_mem[7][70] ), .IN4(n7236), .Q(n4288)
          );
   AO22X1 U3383 (.IN1(n6750), .IN2(n2580), .IN3(\key_mem[8][70] ), .IN4(n6716), .Q(n4289)
          );
   AO22X1 U3384 (.IN1(n7223), .IN2(n2580), .IN3(\key_mem[9][70] ), .IN4(n7213), .Q(n4290)
          );
   AO22X1 U3385 (.IN1(n6797), .IN2(n2580), .IN3(\key_mem[10][70] ), .IN4(n6763), .Q(n4291)
          );
   AO22X1 U3386 (.IN1(n7199), .IN2(n2580), .IN3(\key_mem[11][70] ), .IN4(n7189), .Q(n4292)
          );
   AO22X1 U3387 (.IN1(n6831), .IN2(n2580), .IN3(\key_mem[12][70] ), .IN4(n6841), .Q(n4293)
          );
   AO22X1 U3388 (.IN1(n7178), .IN2(n2580), .IN3(\key_mem[13][70] ), .IN4(n7168), .Q(n4294)
          );
   AO22X1 U3389 (.IN1(n6995), .IN2(n2580), .IN3(\key_mem[14][70] ), .IN4(n7154), .Q(n4295)
          );
   AO221X1 U3390 (.IN1(n7130), .IN2(n2581), .IN3(key[198]), .IN4(n7296), .IN5(n2582), .Q(
          n2580));
   AO222X1 U3391 (.IN1(n7114), .IN2(n2583), .IN3(key[70]), .IN4(n7075), .IN5(n7042), .IN6(
          n2584), .Q(n2582));
   AO22X1 U3392 (.IN1(n7301), .IN2(n2585), .IN3(\key_mem[0][69] ), .IN4(n6933), .Q(n4296)
          );
   AO22X1 U3393 (.IN1(n6809), .IN2(n2585), .IN3(\key_mem[1][69] ), .IN4(n6821), .Q(n4297)
          );
   AO22X1 U3394 (.IN1(n6858), .IN2(n2585), .IN3(\key_mem[2][69] ), .IN4(n6843), .Q(n4298)
          );
   AO22X1 U3395 (.IN1(n6807), .IN2(n2585), .IN3(\key_mem[3][69] ), .IN4(n6863), .Q(n4299)
          );
   AO22X1 U3396 (.IN1(n6888), .IN2(n2585), .IN3(\key_mem[4][69] ), .IN4(n6890), .Q(n4300)
          );
   AO22X1 U3397 (.IN1(n6973), .IN2(n2585), .IN3(\key_mem[5][69] ), .IN4(n7272), .Q(n4301)
          );
   AO22X1 U3398 (.IN1(n7265), .IN2(n2585), .IN3(\key_mem[6][69] ), .IN4(n7258), .Q(n4302)
          );
   AO22X1 U3399 (.IN1(n7246), .IN2(n2585), .IN3(\key_mem[7][69] ), .IN4(n7241), .Q(n4303)
          );
   AO22X1 U3400 (.IN1(n6751), .IN2(n2585), .IN3(\key_mem[8][69] ), .IN4(n6726), .Q(n4304)
          );
   AO22X1 U3401 (.IN1(n6975), .IN2(n2585), .IN3(\key_mem[9][69] ), .IN4(n7216), .Q(n4305)
          );
   AO22X1 U3402 (.IN1(n6798), .IN2(n2585), .IN3(\key_mem[10][69] ), .IN4(n6773), .Q(n4306)
          );
   AO22X1 U3403 (.IN1(n6977), .IN2(n2585), .IN3(\key_mem[11][69] ), .IN4(n7192), .Q(n4307)
          );
   AO22X1 U3404 (.IN1(n6826), .IN2(n2585), .IN3(\key_mem[12][69] ), .IN4(n6984), .Q(n4308)
          );
   AO22X1 U3405 (.IN1(n6979), .IN2(n2585), .IN3(\key_mem[13][69] ), .IN4(n7171), .Q(n4309)
          );
   AO22X1 U3406 (.IN1(n7162), .IN2(n2585), .IN3(\key_mem[14][69] ), .IN4(n7155), .Q(n4310)
          );
   AO221X1 U3407 (.IN1(n7130), .IN2(n2586), .IN3(key[197]), .IN4(n7304), .IN5(n2587), .Q(
          n2585));
   AO222X1 U3408 (.IN1(n7113), .IN2(n2588), .IN3(key[69]), .IN4(n7075), .IN5(n7042), .IN6(
          n2589), .Q(n2587));
   AO22X1 U3409 (.IN1(n7300), .IN2(n2590), .IN3(\key_mem[0][68] ), .IN4(n6933), .Q(n4311)
          );
   AO22X1 U3410 (.IN1(n6927), .IN2(n2590), .IN3(\key_mem[1][68] ), .IN4(n6822), .Q(n4312)
          );
   AO22X1 U3411 (.IN1(n6857), .IN2(n2590), .IN3(\key_mem[2][68] ), .IN4(n6844), .Q(n4313)
          );
   AO22X1 U3412 (.IN1(n6806), .IN2(n2590), .IN3(\key_mem[3][68] ), .IN4(n6861), .Q(n4314)
          );
   AO22X1 U3413 (.IN1(n7288), .IN2(n2590), .IN3(\key_mem[4][68] ), .IN4(n6917), .Q(n4315)
          );
   AO22X1 U3414 (.IN1(n7019), .IN2(n2590), .IN3(\key_mem[5][68] ), .IN4(n7281), .Q(n4316)
          );
   AO22X1 U3415 (.IN1(n7016), .IN2(n2590), .IN3(\key_mem[6][68] ), .IN4(n7259), .Q(n4317)
          );
   AO22X1 U3416 (.IN1(n7247), .IN2(n2590), .IN3(\key_mem[7][68] ), .IN4(n7242), .Q(n4318)
          );
   AO22X1 U3417 (.IN1(n6752), .IN2(n2590), .IN3(\key_mem[8][68] ), .IN4(n6717), .Q(n4319)
          );
   AO22X1 U3418 (.IN1(n7008), .IN2(n2590), .IN3(\key_mem[9][68] ), .IN4(n7225), .Q(n4320)
          );
   AO22X1 U3419 (.IN1(n6799), .IN2(n2590), .IN3(\key_mem[10][68] ), .IN4(n6764), .Q(n4321)
          );
   AO22X1 U3420 (.IN1(n7003), .IN2(n2590), .IN3(\key_mem[11][68] ), .IN4(n7201), .Q(n4322)
          );
   AO22X1 U3421 (.IN1(n6831), .IN2(n2590), .IN3(\key_mem[12][68] ), .IN4(n6839), .Q(n4323)
          );
   AO22X1 U3422 (.IN1(n6998), .IN2(n2590), .IN3(\key_mem[13][68] ), .IN4(n7180), .Q(n4324)
          );
   AO22X1 U3423 (.IN1(n7161), .IN2(n2590), .IN3(\key_mem[14][68] ), .IN4(n7148), .Q(n4325)
          );
   AO221X1 U3424 (.IN1(n7130), .IN2(n2591), .IN3(key[196]), .IN4(n7303), .IN5(n2592), .Q(
          n2590));
   AO222X1 U3425 (.IN1(n7113), .IN2(n2593), .IN3(key[68]), .IN4(n7075), .IN5(n7042), .IN6(
          n2594), .Q(n2592));
   AO22X1 U3426 (.IN1(n7308), .IN2(n2595), .IN3(\key_mem[0][67] ), .IN4(n6933), .Q(n4326)
          );
   AO22X1 U3427 (.IN1(n6808), .IN2(n2595), .IN3(\key_mem[1][67] ), .IN4(n6823), .Q(n4327)
          );
   AO22X1 U3428 (.IN1(n6854), .IN2(n2595), .IN3(\key_mem[2][67] ), .IN4(n6851), .Q(n4328)
          );
   AO22X1 U3429 (.IN1(n6989), .IN2(n2595), .IN3(\key_mem[3][67] ), .IN4(n6867), .Q(n4329)
          );
   AO22X1 U3430 (.IN1(n6916), .IN2(n2595), .IN3(\key_mem[4][67] ), .IN4(n6914), .Q(n4330)
          );
   AO22X1 U3431 (.IN1(n7279), .IN2(n2595), .IN3(\key_mem[5][67] ), .IN4(n7267), .Q(n4331)
          );
   AO22X1 U3432 (.IN1(n7264), .IN2(n2595), .IN3(\key_mem[6][67] ), .IN4(n7258), .Q(n4332)
          );
   AO22X1 U3433 (.IN1(n7248), .IN2(n2595), .IN3(\key_mem[7][67] ), .IN4(n7242), .Q(n4333)
          );
   AO22X1 U3434 (.IN1(n6756), .IN2(n2595), .IN3(\key_mem[8][67] ), .IN4(n6735), .Q(n4334)
          );
   AO22X1 U3435 (.IN1(n7223), .IN2(n2595), .IN3(\key_mem[9][67] ), .IN4(n7211), .Q(n4335)
          );
   AO22X1 U3436 (.IN1(n6803), .IN2(n2595), .IN3(\key_mem[10][67] ), .IN4(n6782), .Q(n4336)
          );
   AO22X1 U3437 (.IN1(n7199), .IN2(n2595), .IN3(\key_mem[11][67] ), .IN4(n7187), .Q(n4337)
          );
   AO22X1 U3438 (.IN1(n6840), .IN2(n2595), .IN3(\key_mem[12][67] ), .IN4(n2289), .Q(n4338)
          );
   AO22X1 U3439 (.IN1(n7178), .IN2(n2595), .IN3(\key_mem[13][67] ), .IN4(n7166), .Q(n4339)
          );
   AO22X1 U3440 (.IN1(n7159), .IN2(n2595), .IN3(\key_mem[14][67] ), .IN4(n7149), .Q(n4340)
          );
   AO221X1 U3441 (.IN1(n7131), .IN2(n2596), .IN3(key[195]), .IN4(n7301), .IN5(n2597), .Q(
          n2595));
   AO222X1 U3442 (.IN1(n7113), .IN2(n2598), .IN3(key[67]), .IN4(n7076), .IN5(n7043), .IN6(
          n2599), .Q(n2597));
   AO22X1 U3443 (.IN1(n7307), .IN2(n2600), .IN3(\key_mem[0][66] ), .IN4(n6933), .Q(n4341)
          );
   AO22X1 U3444 (.IN1(n6927), .IN2(n2600), .IN3(\key_mem[1][66] ), .IN4(n6819), .Q(n4342)
          );
   AO22X1 U3445 (.IN1(n6852), .IN2(n2600), .IN3(\key_mem[2][66] ), .IN4(n6848), .Q(n4343)
          );
   AO22X1 U3446 (.IN1(n6807), .IN2(n2600), .IN3(\key_mem[3][66] ), .IN4(n6868), .Q(n4344)
          );
   AO22X1 U3447 (.IN1(n6922), .IN2(n2600), .IN3(\key_mem[4][66] ), .IN4(n6919), .Q(n4345)
          );
   AO22X1 U3448 (.IN1(n6974), .IN2(n2600), .IN3(\key_mem[5][66] ), .IN4(n7270), .Q(n4346)
          );
   AO22X1 U3449 (.IN1(n7263), .IN2(n2600), .IN3(\key_mem[6][66] ), .IN4(n7255), .Q(n4347)
          );
   AO22X1 U3450 (.IN1(n7250), .IN2(n2600), .IN3(\key_mem[7][66] ), .IN4(n7238), .Q(n4348)
          );
   AO22X1 U3451 (.IN1(n6757), .IN2(n2600), .IN3(\key_mem[8][66] ), .IN4(n6737), .Q(n4349)
          );
   AO22X1 U3452 (.IN1(n6976), .IN2(n2600), .IN3(\key_mem[9][66] ), .IN4(n7213), .Q(n4350)
          );
   AO22X1 U3453 (.IN1(n6804), .IN2(n2600), .IN3(\key_mem[10][66] ), .IN4(n6784), .Q(n4351)
          );
   AO22X1 U3454 (.IN1(n6978), .IN2(n2600), .IN3(\key_mem[11][66] ), .IN4(n7189), .Q(n4352)
          );
   AO22X1 U3455 (.IN1(n6829), .IN2(n2600), .IN3(\key_mem[12][66] ), .IN4(n6984), .Q(n4353)
          );
   AO22X1 U3456 (.IN1(n6980), .IN2(n2600), .IN3(\key_mem[13][66] ), .IN4(n7168), .Q(n4354)
          );
   AO22X1 U3457 (.IN1(n7158), .IN2(n2600), .IN3(\key_mem[14][66] ), .IN4(n7156), .Q(n4355)
          );
   AO221X1 U3458 (.IN1(n7131), .IN2(n2601), .IN3(key[194]), .IN4(n7300), .IN5(n2602), .Q(
          n2600));
   AO222X1 U3459 (.IN1(n7113), .IN2(n2603), .IN3(key[66]), .IN4(n7076), .IN5(n7043), .IN6(
          n2604), .Q(n2602));
   AO22X1 U3460 (.IN1(n7306), .IN2(n2605), .IN3(\key_mem[0][65] ), .IN4(n6933), .Q(n4356)
          );
   AO22X1 U3461 (.IN1(n6810), .IN2(n2605), .IN3(\key_mem[1][65] ), .IN4(n6824), .Q(n4357)
          );
   AO22X1 U3462 (.IN1(n6857), .IN2(n2605), .IN3(\key_mem[2][65] ), .IN4(n6845), .Q(n4358)
          );
   AO22X1 U3463 (.IN1(n6870), .IN2(n2605), .IN3(\key_mem[3][65] ), .IN4(n6860), .Q(n4359)
          );
   AO22X1 U3464 (.IN1(n6921), .IN2(n2605), .IN3(\key_mem[4][65] ), .IN4(n6915), .Q(n4360)
          );
   AO22X1 U3465 (.IN1(n6973), .IN2(n2605), .IN3(\key_mem[5][65] ), .IN4(n2282), .Q(n4361)
          );
   AO22X1 U3466 (.IN1(n7262), .IN2(n2605), .IN3(\key_mem[6][65] ), .IN4(n7257), .Q(n4362)
          );
   AO22X1 U3467 (.IN1(n7249), .IN2(n2605), .IN3(\key_mem[7][65] ), .IN4(n2284), .Q(n4363)
          );
   AO22X1 U3468 (.IN1(n6757), .IN2(n2605), .IN3(\key_mem[8][65] ), .IN4(n6738), .Q(n4364)
          );
   AO22X1 U3469 (.IN1(n6975), .IN2(n2605), .IN3(\key_mem[9][65] ), .IN4(n2286), .Q(n4365)
          );
   AO22X1 U3470 (.IN1(n6804), .IN2(n2605), .IN3(\key_mem[10][65] ), .IN4(n6785), .Q(n4366)
          );
   AO22X1 U3471 (.IN1(n6977), .IN2(n2605), .IN3(\key_mem[11][65] ), .IN4(n2288), .Q(n4367)
          );
   AO22X1 U3472 (.IN1(n6827), .IN2(n2605), .IN3(\key_mem[12][65] ), .IN4(n7185), .Q(n4368)
          );
   AO22X1 U3473 (.IN1(n6979), .IN2(n2605), .IN3(\key_mem[13][65] ), .IN4(n2290), .Q(n4369)
          );
   AO22X1 U3474 (.IN1(n7162), .IN2(n2605), .IN3(\key_mem[14][65] ), .IN4(n7157), .Q(n4370)
          );
   AO221X1 U3475 (.IN1(n7131), .IN2(n2606), .IN3(key[193]), .IN4(n7307), .IN5(n2607), .Q(
          n2605));
   AO222X1 U3476 (.IN1(n7113), .IN2(n2608), .IN3(key[65]), .IN4(n7076), .IN5(n7043), .IN6(
          n2609), .Q(n2607));
   AO22X1 U3477 (.IN1(n7305), .IN2(n2610), .IN3(\key_mem[0][64] ), .IN4(n6933), .Q(n4371)
          );
   AO22X1 U3478 (.IN1(n6811), .IN2(n2610), .IN3(\key_mem[1][64] ), .IN4(n6823), .Q(n4372)
          );
   AO22X1 U3479 (.IN1(n6854), .IN2(n2610), .IN3(\key_mem[2][64] ), .IN4(n6845), .Q(n4373)
          );
   AO22X1 U3480 (.IN1(n6807), .IN2(n2610), .IN3(\key_mem[3][64] ), .IN4(n6861), .Q(n4374)
          );
   AO22X1 U3481 (.IN1(n6924), .IN2(n2610), .IN3(\key_mem[4][64] ), .IN4(n6918), .Q(n4375)
          );
   AO22X1 U3482 (.IN1(n7283), .IN2(n2610), .IN3(\key_mem[5][64] ), .IN4(n7282), .Q(n4376)
          );
   AO22X1 U3483 (.IN1(n7262), .IN2(n2610), .IN3(\key_mem[6][64] ), .IN4(n7254), .Q(n4377)
          );
   AO22X1 U3484 (.IN1(n7247), .IN2(n2610), .IN3(\key_mem[7][64] ), .IN4(n7012), .Q(n4378)
          );
   AO22X1 U3485 (.IN1(n6758), .IN2(n2610), .IN3(\key_mem[8][64] ), .IN4(n6727), .Q(n4379)
          );
   AO22X1 U3486 (.IN1(n7227), .IN2(n2610), .IN3(\key_mem[9][64] ), .IN4(n7226), .Q(n4380)
          );
   AO22X1 U3487 (.IN1(n6805), .IN2(n2610), .IN3(\key_mem[10][64] ), .IN4(n6774), .Q(n4381)
          );
   AO22X1 U3488 (.IN1(n7203), .IN2(n2610), .IN3(\key_mem[11][64] ), .IN4(n7202), .Q(n4382)
          );
   AO22X1 U3489 (.IN1(n6831), .IN2(n2610), .IN3(\key_mem[12][64] ), .IN4(n6841), .Q(n4383)
          );
   AO22X1 U3490 (.IN1(n7182), .IN2(n2610), .IN3(\key_mem[13][64] ), .IN4(n7181), .Q(n4384)
          );
   AO22X1 U3491 (.IN1(n7160), .IN2(n2610), .IN3(\key_mem[14][64] ), .IN4(n7152), .Q(n4385)
          );
   AO221X1 U3492 (.IN1(n7131), .IN2(n2611), .IN3(key[192]), .IN4(n7306), .IN5(n2612), .Q(
          n2610));
   AO222X1 U3493 (.IN1(n7113), .IN2(n2613), .IN3(key[64]), .IN4(n7076), .IN5(n7043), .IN6(
          n2614), .Q(n2612));
   AO22X1 U3494 (.IN1(n7299), .IN2(n2615), .IN3(\key_mem[0][63] ), .IN4(n6933), .Q(n4386)
          );
   AO22X1 U3495 (.IN1(n6810), .IN2(n2615), .IN3(\key_mem[1][63] ), .IN4(n6822), .Q(n4387)
          );
   AO22X1 U3496 (.IN1(n6853), .IN2(n2615), .IN3(\key_mem[2][63] ), .IN4(n6847), .Q(n4388)
          );
   AO22X1 U3497 (.IN1(n6870), .IN2(n2615), .IN3(\key_mem[3][63] ), .IN4(n6876), .Q(n4389)
          );
   AO22X1 U3498 (.IN1(n6889), .IN2(n2615), .IN3(\key_mem[4][63] ), .IN4(n6925), .Q(n4390)
          );
   AO22X1 U3499 (.IN1(n7276), .IN2(n2615), .IN3(\key_mem[5][63] ), .IN4(n7267), .Q(n4391)
          );
   AO22X1 U3500 (.IN1(n7262), .IN2(n2615), .IN3(\key_mem[6][63] ), .IN4(n7259), .Q(n4392)
          );
   AO22X1 U3501 (.IN1(n7247), .IN2(n2615), .IN3(\key_mem[7][63] ), .IN4(n7243), .Q(n4393)
          );
   AO22X1 U3502 (.IN1(n6748), .IN2(n2615), .IN3(\key_mem[8][63] ), .IN4(n6725), .Q(n4394)
          );
   AO22X1 U3503 (.IN1(n7220), .IN2(n2615), .IN3(\key_mem[9][63] ), .IN4(n7211), .Q(n4395)
          );
   AO22X1 U3504 (.IN1(n6795), .IN2(n2615), .IN3(\key_mem[10][63] ), .IN4(n6772), .Q(n4396)
          );
   AO22X1 U3505 (.IN1(n7196), .IN2(n2615), .IN3(\key_mem[11][63] ), .IN4(n7187), .Q(n4397)
          );
   AO22X1 U3506 (.IN1(n6829), .IN2(n2615), .IN3(\key_mem[12][63] ), .IN4(n6833), .Q(n4398)
          );
   AO22X1 U3507 (.IN1(n7175), .IN2(n2615), .IN3(\key_mem[13][63] ), .IN4(n7166), .Q(n4399)
          );
   AO22X1 U3508 (.IN1(n7161), .IN2(n2615), .IN3(\key_mem[14][63] ), .IN4(n7157), .Q(n4400)
          );
   AO221X1 U3509 (.IN1(n7131), .IN2(n2616), .IN3(key[191]), .IN4(n7292), .IN5(n2617), .Q(
          n2615));
   AO222X1 U3510 (.IN1(n7113), .IN2(n2618), .IN3(key[63]), .IN4(n7076), .IN5(n7043), .IN6(
          n2619), .Q(n2617));
   AO22X1 U3511 (.IN1(n7298), .IN2(n2620), .IN3(\key_mem[0][62] ), .IN4(n6933), .Q(n4401)
          );
   AO22X1 U3512 (.IN1(n6811), .IN2(n2620), .IN3(\key_mem[1][62] ), .IN4(n6824), .Q(n4402)
          );
   AO22X1 U3513 (.IN1(n6858), .IN2(n2620), .IN3(\key_mem[2][62] ), .IN4(n6842), .Q(n4403)
          );
   AO22X1 U3514 (.IN1(n6989), .IN2(n2620), .IN3(\key_mem[3][62] ), .IN4(n6863), .Q(n4404)
          );
   AO22X1 U3515 (.IN1(n7022), .IN2(n2620), .IN3(\key_mem[4][62] ), .IN4(n7284), .Q(n4405)
          );
   AO22X1 U3516 (.IN1(n7020), .IN2(n2620), .IN3(\key_mem[5][62] ), .IN4(n7269), .Q(n4406)
          );
   AO22X1 U3517 (.IN1(n7017), .IN2(n2620), .IN3(\key_mem[6][62] ), .IN4(n7258), .Q(n4407)
          );
   AO22X1 U3518 (.IN1(n7244), .IN2(n2620), .IN3(\key_mem[7][62] ), .IN4(n7235), .Q(n4408)
          );
   AO22X1 U3519 (.IN1(n6749), .IN2(n2620), .IN3(\key_mem[8][62] ), .IN4(n6724), .Q(n4409)
          );
   AO22X1 U3520 (.IN1(n7009), .IN2(n2620), .IN3(\key_mem[9][62] ), .IN4(n7212), .Q(n4410)
          );
   AO22X1 U3521 (.IN1(n6796), .IN2(n2620), .IN3(\key_mem[10][62] ), .IN4(n6771), .Q(n4411)
          );
   AO22X1 U3522 (.IN1(n7004), .IN2(n2620), .IN3(\key_mem[11][62] ), .IN4(n7188), .Q(n4412)
          );
   AO22X1 U3523 (.IN1(n6987), .IN2(n2620), .IN3(\key_mem[12][62] ), .IN4(n6983), .Q(n4413)
          );
   AO22X1 U3524 (.IN1(n6999), .IN2(n2620), .IN3(\key_mem[13][62] ), .IN4(n7167), .Q(n4414)
          );
   AO22X1 U3525 (.IN1(n7164), .IN2(n2620), .IN3(\key_mem[14][62] ), .IN4(n7165), .Q(n4415)
          );
   AO221X1 U3526 (.IN1(n7131), .IN2(n2621), .IN3(key[190]), .IN4(n7297), .IN5(n2622), .Q(
          n2620));
   AO222X1 U3527 (.IN1(n7113), .IN2(n2623), .IN3(key[62]), .IN4(n7076), .IN5(n7043), .IN6(
          n2624), .Q(n2622));
   AO22X1 U3528 (.IN1(n7297), .IN2(n2625), .IN3(\key_mem[0][61] ), .IN4(n6933), .Q(n4416)
          );
   AO22X1 U3529 (.IN1(n6926), .IN2(n2625), .IN3(\key_mem[1][61] ), .IN4(n6824), .Q(n4417)
          );
   AO22X1 U3530 (.IN1(n6853), .IN2(n2625), .IN3(\key_mem[2][61] ), .IN4(n6849), .Q(n4418)
          );
   AO22X1 U3531 (.IN1(n6807), .IN2(n2625), .IN3(\key_mem[3][61] ), .IN4(n6863), .Q(n4419)
          );
   AO22X1 U3532 (.IN1(n6990), .IN2(n2625), .IN3(\key_mem[4][61] ), .IN4(n7021), .Q(n4420)
          );
   AO22X1 U3533 (.IN1(n7278), .IN2(n2625), .IN3(\key_mem[5][61] ), .IN4(n2282), .Q(n4421)
          );
   AO22X1 U3534 (.IN1(n6970), .IN2(n2625), .IN3(\key_mem[6][61] ), .IN4(n7256), .Q(n4422)
          );
   AO22X1 U3535 (.IN1(n7248), .IN2(n2625), .IN3(\key_mem[7][61] ), .IN4(n7236), .Q(n4423)
          );
   AO22X1 U3536 (.IN1(n6750), .IN2(n2625), .IN3(\key_mem[8][61] ), .IN4(n6721), .Q(n4424)
          );
   AO22X1 U3537 (.IN1(n7222), .IN2(n2625), .IN3(\key_mem[9][61] ), .IN4(n2286), .Q(n4425)
          );
   AO22X1 U3538 (.IN1(n6797), .IN2(n2625), .IN3(\key_mem[10][61] ), .IN4(n6768), .Q(n4426)
          );
   AO22X1 U3539 (.IN1(n7198), .IN2(n2625), .IN3(\key_mem[11][61] ), .IN4(n2288), .Q(n4427)
          );
   AO22X1 U3540 (.IN1(n7183), .IN2(n2625), .IN3(\key_mem[12][61] ), .IN4(n6838), .Q(n4428)
          );
   AO22X1 U3541 (.IN1(n7177), .IN2(n2625), .IN3(\key_mem[13][61] ), .IN4(n2290), .Q(n4429)
          );
   AO22X1 U3542 (.IN1(n7163), .IN2(n2625), .IN3(\key_mem[14][61] ), .IN4(n7150), .Q(n4430)
          );
   AO222X1 U3544 (.IN1(n7113), .IN2(n2628), .IN3(key[61]), .IN4(n7076), .IN5(n7043), .IN6(
          n2629), .Q(n2627));
   AO22X1 U3545 (.IN1(n7296), .IN2(n2630), .IN3(\key_mem[0][60] ), .IN4(n6933), .Q(n4431)
          );
   AO22X1 U3546 (.IN1(n6808), .IN2(n2630), .IN3(\key_mem[1][60] ), .IN4(n6825), .Q(n4432)
          );
   AO22X1 U3547 (.IN1(n6855), .IN2(n2630), .IN3(\key_mem[2][60] ), .IN4(n6846), .Q(n4433)
          );
   AO22X1 U3548 (.IN1(n6870), .IN2(n2630), .IN3(\key_mem[3][60] ), .IN4(n6862), .Q(n4434)
          );
   AO22X1 U3549 (.IN1(n6889), .IN2(n2630), .IN3(\key_mem[4][60] ), .IN4(n6923), .Q(n4435)
          );
   AO22X1 U3550 (.IN1(n6974), .IN2(n2630), .IN3(\key_mem[5][60] ), .IN4(n7282), .Q(n4436)
          );
   AO22X1 U3551 (.IN1(n6969), .IN2(n2630), .IN3(\key_mem[6][60] ), .IN4(n7257), .Q(n4437)
          );
   AO22X1 U3552 (.IN1(n7013), .IN2(n2630), .IN3(\key_mem[7][60] ), .IN4(n7240), .Q(n4438)
          );
   AO22X1 U3553 (.IN1(n6754), .IN2(n2630), .IN3(\key_mem[8][60] ), .IN4(n6722), .Q(n4439)
          );
   AO22X1 U3554 (.IN1(n6976), .IN2(n2630), .IN3(\key_mem[9][60] ), .IN4(n7226), .Q(n4440)
          );
   AO22X1 U3555 (.IN1(n6801), .IN2(n2630), .IN3(\key_mem[10][60] ), .IN4(n6769), .Q(n4441)
          );
   AO22X1 U3556 (.IN1(n6978), .IN2(n2630), .IN3(\key_mem[11][60] ), .IN4(n7202), .Q(n4442)
          );
   AO22X1 U3557 (.IN1(n6840), .IN2(n2630), .IN3(\key_mem[12][60] ), .IN4(n6839), .Q(n4443)
          );
   AO22X1 U3558 (.IN1(n6980), .IN2(n2630), .IN3(\key_mem[13][60] ), .IN4(n7181), .Q(n4444)
          );
   AO22X1 U3559 (.IN1(n6972), .IN2(n2630), .IN3(\key_mem[14][60] ), .IN4(n7147), .Q(n4445)
          );
   AO222X1 U3561 (.IN1(n7113), .IN2(n2633), .IN3(key[60]), .IN4(n7076), .IN5(n7043), .IN6(
          n2634), .Q(n2632));
   AO22X1 U3562 (.IN1(n7295), .IN2(n2635), .IN3(\key_mem[0][59] ), .IN4(n6932), .Q(n4446)
          );
   AO22X1 U3563 (.IN1(n6811), .IN2(n2635), .IN3(\key_mem[1][59] ), .IN4(n6822), .Q(n4447)
          );
   AO22X1 U3564 (.IN1(n6856), .IN2(n2635), .IN3(\key_mem[2][59] ), .IN4(n6843), .Q(n4448)
          );
   AO22X1 U3565 (.IN1(n6873), .IN2(n2635), .IN3(\key_mem[3][59] ), .IN4(n6864), .Q(n4449)
          );
   AO22X1 U3566 (.IN1(n6922), .IN2(n2635), .IN3(\key_mem[4][59] ), .IN4(n6919), .Q(n4450)
          );
   AO22X1 U3567 (.IN1(n7277), .IN2(n2635), .IN3(\key_mem[5][59] ), .IN4(n7271), .Q(n4451)
          );
   AO22X1 U3568 (.IN1(n7016), .IN2(n2635), .IN3(\key_mem[6][59] ), .IN4(n7256), .Q(n4452)
          );
   AO22X1 U3569 (.IN1(n7014), .IN2(n2635), .IN3(\key_mem[7][59] ), .IN4(n7236), .Q(n4453)
          );
   AO22X1 U3570 (.IN1(n6755), .IN2(n2635), .IN3(\key_mem[8][59] ), .IN4(n6742), .Q(n4454)
          );
   AO22X1 U3571 (.IN1(n7221), .IN2(n2635), .IN3(\key_mem[9][59] ), .IN4(n7215), .Q(n4455)
          );
   AO22X1 U3572 (.IN1(n6802), .IN2(n2635), .IN3(\key_mem[10][59] ), .IN4(n6789), .Q(n4456)
          );
   AO22X1 U3573 (.IN1(n7197), .IN2(n2635), .IN3(\key_mem[11][59] ), .IN4(n7191), .Q(n4457)
          );
   AO22X1 U3574 (.IN1(n7186), .IN2(n2635), .IN3(\key_mem[12][59] ), .IN4(n6834), .Q(n4458)
          );
   AO22X1 U3575 (.IN1(n7176), .IN2(n2635), .IN3(\key_mem[13][59] ), .IN4(n7170), .Q(n4459)
          );
   AO22X1 U3576 (.IN1(n7164), .IN2(n2635), .IN3(\key_mem[14][59] ), .IN4(n7165), .Q(n4460)
          );
   AO221X1 U3577 (.IN1(n7131), .IN2(n2636), .IN3(key[187]), .IN4(n7306), .IN5(n2637), .Q(
          n2635));
   AO222X1 U3578 (.IN1(n7113), .IN2(n2638), .IN3(key[59]), .IN4(n7076), .IN5(n7043), .IN6(
          n2639), .Q(n2637));
   AO22X1 U3579 (.IN1(n7304), .IN2(n2640), .IN3(\key_mem[0][58] ), .IN4(n6932), .Q(n4461)
          );
   AO22X1 U3580 (.IN1(n6813), .IN2(n2640), .IN3(\key_mem[1][58] ), .IN4(n6818), .Q(n4462)
          );
   AO22X1 U3581 (.IN1(n6988), .IN2(n2640), .IN3(\key_mem[2][58] ), .IN4(n6842), .Q(n4463)
          );
   AO22X1 U3582 (.IN1(n6869), .IN2(n2640), .IN3(\key_mem[3][58] ), .IN4(n6860), .Q(n4464)
          );
   AO22X1 U3583 (.IN1(n6924), .IN2(n2640), .IN3(\key_mem[4][58] ), .IN4(n6915), .Q(n4465)
          );
   AO22X1 U3584 (.IN1(n6974), .IN2(n2640), .IN3(\key_mem[5][58] ), .IN4(n7272), .Q(n4466)
          );
   AO22X1 U3585 (.IN1(n7017), .IN2(n2640), .IN3(\key_mem[6][58] ), .IN4(n7015), .Q(n4467)
          );
   AO22X1 U3586 (.IN1(n7244), .IN2(n2640), .IN3(\key_mem[7][58] ), .IN4(n7243), .Q(n4468)
          );
   AO22X1 U3587 (.IN1(n6756), .IN2(n2640), .IN3(\key_mem[8][58] ), .IN4(n6727), .Q(n4469)
          );
   AO22X1 U3588 (.IN1(n6976), .IN2(n2640), .IN3(\key_mem[9][58] ), .IN4(n7216), .Q(n4470)
          );
   AO22X1 U3589 (.IN1(n6803), .IN2(n2640), .IN3(\key_mem[10][58] ), .IN4(n6774), .Q(n4471)
          );
   AO22X1 U3590 (.IN1(n6978), .IN2(n2640), .IN3(\key_mem[11][58] ), .IN4(n7192), .Q(n4472)
          );
   AO22X1 U3591 (.IN1(n6835), .IN2(n2640), .IN3(\key_mem[12][58] ), .IN4(n6982), .Q(n4473)
          );
   AO22X1 U3592 (.IN1(n6980), .IN2(n2640), .IN3(\key_mem[13][58] ), .IN4(n7171), .Q(n4474)
          );
   AO22X1 U3593 (.IN1(n6996), .IN2(n2640), .IN3(\key_mem[14][58] ), .IN4(n6994), .Q(n4475)
          );
   AO222X1 U3595 (.IN1(n7113), .IN2(n2643), .IN3(key[58]), .IN4(n7076), .IN5(n7043), .IN6(
          n2644), .Q(n2642));
   AO22X1 U3596 (.IN1(n7303), .IN2(n2645), .IN3(\key_mem[0][57] ), .IN4(n6932), .Q(n4476)
          );
   AO22X1 U3597 (.IN1(n6810), .IN2(n2645), .IN3(\key_mem[1][57] ), .IN4(n6823), .Q(n4477)
          );
   AO22X1 U3598 (.IN1(n6856), .IN2(n2645), .IN3(\key_mem[2][57] ), .IN4(n6846), .Q(n4478)
          );
   AO22X1 U3599 (.IN1(n6806), .IN2(n2645), .IN3(\key_mem[3][57] ), .IN4(n6866), .Q(n4479)
          );
   AO22X1 U3600 (.IN1(n6888), .IN2(n2645), .IN3(\key_mem[4][57] ), .IN4(n6915), .Q(n4480)
          );
   AO22X1 U3601 (.IN1(n7283), .IN2(n2645), .IN3(\key_mem[5][57] ), .IN4(n7282), .Q(n4481)
          );
   AO22X1 U3602 (.IN1(n7017), .IN2(n2645), .IN3(\key_mem[6][57] ), .IN4(n7251), .Q(n4482)
          );
   AO22X1 U3603 (.IN1(n7245), .IN2(n2645), .IN3(\key_mem[7][57] ), .IN4(n7237), .Q(n4483)
          );
   AO22X1 U3604 (.IN1(n6758), .IN2(n2645), .IN3(\key_mem[8][57] ), .IN4(n6729), .Q(n4484)
          );
   AO22X1 U3605 (.IN1(n7227), .IN2(n2645), .IN3(\key_mem[9][57] ), .IN4(n7226), .Q(n4485)
          );
   AO22X1 U3606 (.IN1(n6805), .IN2(n2645), .IN3(\key_mem[10][57] ), .IN4(n6776), .Q(n4486)
          );
   AO22X1 U3607 (.IN1(n7203), .IN2(n2645), .IN3(\key_mem[11][57] ), .IN4(n7202), .Q(n4487)
          );
   AO22X1 U3608 (.IN1(n6826), .IN2(n2645), .IN3(\key_mem[12][57] ), .IN4(n6828), .Q(n4488)
          );
   AO22X1 U3609 (.IN1(n7182), .IN2(n2645), .IN3(\key_mem[13][57] ), .IN4(n7181), .Q(n4489)
          );
   AO22X1 U3610 (.IN1(n7160), .IN2(n2645), .IN3(\key_mem[14][57] ), .IN4(n7149), .Q(n4490)
          );
   AO222X1 U3612 (.IN1(n7113), .IN2(n2648), .IN3(key[57]), .IN4(n7076), .IN5(n7043), .IN6(
          n2649), .Q(n2647));
   AO22X1 U3613 (.IN1(n7302), .IN2(n2650), .IN3(\key_mem[0][56] ), .IN4(n6932), .Q(n4491)
          );
   AO22X1 U3614 (.IN1(n6809), .IN2(n2650), .IN3(\key_mem[1][56] ), .IN4(n6819), .Q(n4492)
          );
   AO22X1 U3615 (.IN1(n6854), .IN2(n2650), .IN3(\key_mem[2][56] ), .IN4(n6845), .Q(n4493)
          );
   AO22X1 U3616 (.IN1(n6875), .IN2(n2650), .IN3(\key_mem[3][56] ), .IN4(n6876), .Q(n4494)
          );
   AO22X1 U3617 (.IN1(n6922), .IN2(n2650), .IN3(\key_mem[4][56] ), .IN4(n6917), .Q(n4495)
          );
   AO22X1 U3618 (.IN1(n7020), .IN2(n2650), .IN3(\key_mem[5][56] ), .IN4(n2282), .Q(n4496)
          );
   AO22X1 U3619 (.IN1(n7262), .IN2(n2650), .IN3(\key_mem[6][56] ), .IN4(n7256), .Q(n4497)
          );
   AO22X1 U3620 (.IN1(n7246), .IN2(n2650), .IN3(\key_mem[7][56] ), .IN4(n7237), .Q(n4498)
          );
   AO22X1 U3621 (.IN1(n6748), .IN2(n2650), .IN3(\key_mem[8][56] ), .IN4(n6730), .Q(n4499)
          );
   AO22X1 U3622 (.IN1(n7009), .IN2(n2650), .IN3(\key_mem[9][56] ), .IN4(n2286), .Q(n4500)
          );
   AO22X1 U3623 (.IN1(n6795), .IN2(n2650), .IN3(\key_mem[10][56] ), .IN4(n6777), .Q(n4501)
          );
   AO22X1 U3624 (.IN1(n7004), .IN2(n2650), .IN3(\key_mem[11][56] ), .IN4(n2288), .Q(n4502)
          );
   AO22X1 U3625 (.IN1(n6832), .IN2(n2650), .IN3(\key_mem[12][56] ), .IN4(n6983), .Q(n4503)
          );
   AO22X1 U3626 (.IN1(n6999), .IN2(n2650), .IN3(\key_mem[13][56] ), .IN4(n2290), .Q(n4504)
          );
   AO22X1 U3627 (.IN1(n7164), .IN2(n2650), .IN3(\key_mem[14][56] ), .IN4(n6994), .Q(n4505)
          );
   AO222X1 U3629 (.IN1(n7112), .IN2(n2653), .IN3(key[56]), .IN4(n7076), .IN5(n7043), .IN6(
          n2654), .Q(n2652));
   AO22X1 U3630 (.IN1(n7301), .IN2(n2655), .IN3(\key_mem[0][55] ), .IN4(n6932), .Q(n4506)
          );
   AO22X1 U3631 (.IN1(n6812), .IN2(n2655), .IN3(\key_mem[1][55] ), .IN4(n6824), .Q(n4507)
          );
   AO22X1 U3632 (.IN1(n6855), .IN2(n2655), .IN3(\key_mem[2][55] ), .IN4(n6847), .Q(n4508)
          );
   AO22X1 U3633 (.IN1(n6873), .IN2(n2655), .IN3(\key_mem[3][55] ), .IN4(n6868), .Q(n4509)
          );
   AO22X1 U3634 (.IN1(n6886), .IN2(n2655), .IN3(\key_mem[4][55] ), .IN4(n6914), .Q(n4510)
          );
   AO22X1 U3635 (.IN1(n6973), .IN2(n2655), .IN3(\key_mem[5][55] ), .IN4(n7269), .Q(n4511)
          );
   AO22X1 U3636 (.IN1(n7261), .IN2(n2655), .IN3(\key_mem[6][55] ), .IN4(n7015), .Q(n4512)
          );
   AO22X1 U3637 (.IN1(n7248), .IN2(n2655), .IN3(\key_mem[7][55] ), .IN4(n7238), .Q(n4513)
          );
   AO22X1 U3638 (.IN1(n6751), .IN2(n2655), .IN3(\key_mem[8][55] ), .IN4(n6717), .Q(n4514)
          );
   AO22X1 U3639 (.IN1(n6975), .IN2(n2655), .IN3(\key_mem[9][55] ), .IN4(n7214), .Q(n4515)
          );
   AO22X1 U3640 (.IN1(n6798), .IN2(n2655), .IN3(\key_mem[10][55] ), .IN4(n6764), .Q(n4516)
          );
   AO22X1 U3641 (.IN1(n6977), .IN2(n2655), .IN3(\key_mem[11][55] ), .IN4(n7190), .Q(n4517)
          );
   AO22X1 U3642 (.IN1(n6987), .IN2(n2655), .IN3(\key_mem[12][55] ), .IN4(n6830), .Q(n4518)
          );
   AO22X1 U3643 (.IN1(n6979), .IN2(n2655), .IN3(\key_mem[13][55] ), .IN4(n7169), .Q(n4519)
          );
   AO22X1 U3644 (.IN1(n7161), .IN2(n2655), .IN3(\key_mem[14][55] ), .IN4(n7149), .Q(n4520)
          );
   AO221X1 U3645 (.IN1(n7132), .IN2(n2656), .IN3(key[183]), .IN4(n2276), .IN5(n2657), .Q(
          n2655));
   AO222X1 U3646 (.IN1(n7112), .IN2(n2658), .IN3(key[55]), .IN4(n7077), .IN5(n7044), .IN6(
          n2659), .Q(n2657));
   AO22X1 U3647 (.IN1(n7300), .IN2(n2660), .IN3(\key_mem[0][54] ), .IN4(n6932), .Q(n4521)
          );
   AO22X1 U3648 (.IN1(n6810), .IN2(n2660), .IN3(\key_mem[1][54] ), .IN4(n6824), .Q(n4522)
          );
   AO22X1 U3649 (.IN1(n6856), .IN2(n2660), .IN3(\key_mem[2][54] ), .IN4(n6843), .Q(n4523)
          );
   AO22X1 U3650 (.IN1(n6869), .IN2(n2660), .IN3(\key_mem[3][54] ), .IN4(n6877), .Q(n4524)
          );
   AO22X1 U3651 (.IN1(n7287), .IN2(n2660), .IN3(\key_mem[4][54] ), .IN4(n6917), .Q(n4525)
          );
   AO22X1 U3652 (.IN1(n7283), .IN2(n2660), .IN3(\key_mem[5][54] ), .IN4(n7271), .Q(n4526)
          );
   AO22X1 U3653 (.IN1(n7261), .IN2(n2660), .IN3(\key_mem[6][54] ), .IN4(n7253), .Q(n4527)
          );
   AO22X1 U3654 (.IN1(n7248), .IN2(n2660), .IN3(\key_mem[7][54] ), .IN4(n7239), .Q(n4528)
          );
   AO22X1 U3655 (.IN1(n6752), .IN2(n2660), .IN3(\key_mem[8][54] ), .IN4(n6718), .Q(n4529)
          );
   AO22X1 U3656 (.IN1(n7227), .IN2(n2660), .IN3(\key_mem[9][54] ), .IN4(n7215), .Q(n4530)
          );
   AO22X1 U3657 (.IN1(n6799), .IN2(n2660), .IN3(\key_mem[10][54] ), .IN4(n6765), .Q(n4531)
          );
   AO22X1 U3658 (.IN1(n7203), .IN2(n2660), .IN3(\key_mem[11][54] ), .IN4(n7191), .Q(n4532)
          );
   AO22X1 U3659 (.IN1(n6840), .IN2(n2660), .IN3(\key_mem[12][54] ), .IN4(n7000), .Q(n4533)
          );
   AO22X1 U3660 (.IN1(n7182), .IN2(n2660), .IN3(\key_mem[13][54] ), .IN4(n7170), .Q(n4534)
          );
   AO22X1 U3661 (.IN1(n7160), .IN2(n2660), .IN3(\key_mem[14][54] ), .IN4(n7155), .Q(n4535)
          );
   AO221X1 U3662 (.IN1(n7132), .IN2(n2661), .IN3(key[182]), .IN4(n7305), .IN5(n2662), .Q(
          n2660));
   AO222X1 U3663 (.IN1(n7112), .IN2(n2663), .IN3(key[54]), .IN4(n7077), .IN5(n7044), .IN6(
          n2664), .Q(n2662));
   AO22X1 U3664 (.IN1(n7304), .IN2(n2665), .IN3(\key_mem[0][53] ), .IN4(n6932), .Q(n4536)
          );
   AO22X1 U3665 (.IN1(n6811), .IN2(n2665), .IN3(\key_mem[1][53] ), .IN4(n6817), .Q(n4537)
          );
   AO22X1 U3666 (.IN1(n6858), .IN2(n2665), .IN3(\key_mem[2][53] ), .IN4(n6859), .Q(n4538)
          );
   AO22X1 U3667 (.IN1(n6806), .IN2(n2665), .IN3(\key_mem[3][53] ), .IN4(n6863), .Q(n4539)
          );
   AO22X1 U3668 (.IN1(n6889), .IN2(n2665), .IN3(\key_mem[4][53] ), .IN4(n6917), .Q(n4540)
          );
   AO22X1 U3669 (.IN1(n7019), .IN2(n2665), .IN3(\key_mem[5][53] ), .IN4(n7018), .Q(n4541)
          );
   AO22X1 U3670 (.IN1(n7261), .IN2(n2665), .IN3(\key_mem[6][53] ), .IN4(n7252), .Q(n4542)
          );
   AO22X1 U3671 (.IN1(n7245), .IN2(n2665), .IN3(\key_mem[7][53] ), .IN4(n7240), .Q(n4543)
          );
   AO22X1 U3672 (.IN1(n6754), .IN2(n2665), .IN3(\key_mem[8][53] ), .IN4(n6719), .Q(n4544)
          );
   AO22X1 U3673 (.IN1(n7008), .IN2(n2665), .IN3(\key_mem[9][53] ), .IN4(n7007), .Q(n4545)
          );
   AO22X1 U3674 (.IN1(n6801), .IN2(n2665), .IN3(\key_mem[10][53] ), .IN4(n6766), .Q(n4546)
          );
   AO22X1 U3675 (.IN1(n7003), .IN2(n2665), .IN3(\key_mem[11][53] ), .IN4(n7002), .Q(n4547)
          );
   AO22X1 U3676 (.IN1(n7183), .IN2(n2665), .IN3(\key_mem[12][53] ), .IN4(n6830), .Q(n4548)
          );
   AO22X1 U3677 (.IN1(n6998), .IN2(n2665), .IN3(\key_mem[13][53] ), .IN4(n6997), .Q(n4549)
          );
   AO22X1 U3678 (.IN1(n7164), .IN2(n2665), .IN3(\key_mem[14][53] ), .IN4(n7152), .Q(n4550)
          );
   AO221X1 U3679 (.IN1(n7132), .IN2(n2666), .IN3(key[181]), .IN4(n7311), .IN5(n2667), .Q(
          n2665));
   AO222X1 U3680 (.IN1(n7112), .IN2(n2668), .IN3(key[53]), .IN4(n7077), .IN5(n7044), .IN6(
          n2669), .Q(n2667));
   AO22X1 U3681 (.IN1(n7303), .IN2(n2670), .IN3(\key_mem[0][52] ), .IN4(n6932), .Q(n4551)
          );
   AO22X1 U3682 (.IN1(n6811), .IN2(n2670), .IN3(\key_mem[1][52] ), .IN4(n6820), .Q(n4552)
          );
   AO22X1 U3683 (.IN1(n6858), .IN2(n2670), .IN3(\key_mem[2][52] ), .IN4(n6850), .Q(n4553)
          );
   AO22X1 U3684 (.IN1(n6869), .IN2(n2670), .IN3(\key_mem[3][52] ), .IN4(n6860), .Q(n4554)
          );
   AO22X1 U3685 (.IN1(n6921), .IN2(n2670), .IN3(\key_mem[4][52] ), .IN4(n6925), .Q(n4555)
          );
   AO22X1 U3686 (.IN1(n7020), .IN2(n2670), .IN3(\key_mem[5][52] ), .IN4(n7281), .Q(n4556)
          );
   AO22X1 U3687 (.IN1(n7261), .IN2(n2670), .IN3(\key_mem[6][52] ), .IN4(n7253), .Q(n4557)
          );
   AO22X1 U3688 (.IN1(n7250), .IN2(n2670), .IN3(\key_mem[7][52] ), .IN4(n7241), .Q(n4558)
          );
   AO22X1 U3689 (.IN1(n6755), .IN2(n2670), .IN3(\key_mem[8][52] ), .IN4(n6720), .Q(n4559)
          );
   AO22X1 U3690 (.IN1(n7009), .IN2(n2670), .IN3(\key_mem[9][52] ), .IN4(n7225), .Q(n4560)
          );
   AO22X1 U3691 (.IN1(n6802), .IN2(n2670), .IN3(\key_mem[10][52] ), .IN4(n6767), .Q(n4561)
          );
   AO22X1 U3692 (.IN1(n7004), .IN2(n2670), .IN3(\key_mem[11][52] ), .IN4(n7201), .Q(n4562)
          );
   AO22X1 U3693 (.IN1(n7001), .IN2(n2670), .IN3(\key_mem[12][52] ), .IN4(n6830), .Q(n4563)
          );
   AO22X1 U3694 (.IN1(n6999), .IN2(n2670), .IN3(\key_mem[13][52] ), .IN4(n7180), .Q(n4564)
          );
   AO22X1 U3695 (.IN1(n6972), .IN2(n2670), .IN3(\key_mem[14][52] ), .IN4(n6994), .Q(n4565)
          );
   AO221X1 U3696 (.IN1(n7132), .IN2(n2671), .IN3(key[180]), .IN4(n7312), .IN5(n2672), .Q(
          n2670));
   AO222X1 U3697 (.IN1(n7112), .IN2(n2673), .IN3(key[52]), .IN4(n7077), .IN5(n7044), .IN6(
          n2674), .Q(n2672));
   AO22X1 U3698 (.IN1(n7302), .IN2(n2675), .IN3(\key_mem[0][51] ), .IN4(n6932), .Q(n4566)
          );
   AO22X1 U3699 (.IN1(n6926), .IN2(n2675), .IN3(\key_mem[1][51] ), .IN4(n6819), .Q(n4567)
          );
   AO22X1 U3700 (.IN1(n6852), .IN2(n2675), .IN3(\key_mem[2][51] ), .IN4(n6848), .Q(n4568)
          );
   AO22X1 U3701 (.IN1(n6806), .IN2(n2675), .IN3(\key_mem[3][51] ), .IN4(n6860), .Q(n4569)
          );
   AO22X1 U3702 (.IN1(n7288), .IN2(n2675), .IN3(\key_mem[4][51] ), .IN4(n6890), .Q(n4570)
          );
   AO22X1 U3703 (.IN1(n7277), .IN2(n2675), .IN3(\key_mem[5][51] ), .IN4(n7018), .Q(n4571)
          );
   AO22X1 U3704 (.IN1(n7266), .IN2(n2675), .IN3(\key_mem[6][51] ), .IN4(n7256), .Q(n4572)
          );
   AO22X1 U3705 (.IN1(n7247), .IN2(n2675), .IN3(\key_mem[7][51] ), .IN4(n7242), .Q(n4573)
          );
   AO22X1 U3706 (.IN1(n6756), .IN2(n2675), .IN3(\key_mem[8][51] ), .IN4(n6721), .Q(n4574)
          );
   AO22X1 U3707 (.IN1(n7221), .IN2(n2675), .IN3(\key_mem[9][51] ), .IN4(n7007), .Q(n4575)
          );
   AO22X1 U3708 (.IN1(n6803), .IN2(n2675), .IN3(\key_mem[10][51] ), .IN4(n6768), .Q(n4576)
          );
   AO22X1 U3709 (.IN1(n7197), .IN2(n2675), .IN3(\key_mem[11][51] ), .IN4(n7002), .Q(n4577)
          );
   AO22X1 U3710 (.IN1(n6835), .IN2(n2675), .IN3(\key_mem[12][51] ), .IN4(n6830), .Q(n4578)
          );
   AO22X1 U3711 (.IN1(n7176), .IN2(n2675), .IN3(\key_mem[13][51] ), .IN4(n6997), .Q(n4579)
          );
   AO22X1 U3712 (.IN1(n7160), .IN2(n2675), .IN3(\key_mem[14][51] ), .IN4(n7150), .Q(n4580)
          );
   AO221X1 U3713 (.IN1(n7132), .IN2(n2676), .IN3(key[179]), .IN4(n7294), .IN5(n2677), .Q(
          n2675));
   AO222X1 U3714 (.IN1(n7112), .IN2(n2678), .IN3(key[51]), .IN4(n7077), .IN5(n7044), .IN6(
          n2679), .Q(n2677));
   AO22X1 U3715 (.IN1(n7301), .IN2(n2680), .IN3(\key_mem[0][50] ), .IN4(n6932), .Q(n4581)
          );
   AO22X1 U3716 (.IN1(n6927), .IN2(n2680), .IN3(\key_mem[1][50] ), .IN4(n6824), .Q(n4582)
          );
   AO22X1 U3717 (.IN1(n6853), .IN2(n2680), .IN3(\key_mem[2][50] ), .IN4(n6850), .Q(n4583)
          );
   AO22X1 U3718 (.IN1(n6873), .IN2(n2680), .IN3(\key_mem[3][50] ), .IN4(n6862), .Q(n4584)
          );
   AO22X1 U3719 (.IN1(n6889), .IN2(n2680), .IN3(\key_mem[4][50] ), .IN4(n6923), .Q(n4585)
          );
   AO22X1 U3720 (.IN1(n7280), .IN2(n2680), .IN3(\key_mem[5][50] ), .IN4(n7267), .Q(n4586)
          );
   AO22X1 U3721 (.IN1(n7266), .IN2(n2680), .IN3(\key_mem[6][50] ), .IN4(n2283), .Q(n4587)
          );
   AO22X1 U3722 (.IN1(n7248), .IN2(n2680), .IN3(\key_mem[7][50] ), .IN4(n7243), .Q(n4588)
          );
   AO22X1 U3723 (.IN1(n6757), .IN2(n2680), .IN3(\key_mem[8][50] ), .IN4(n6726), .Q(n4589)
          );
   AO22X1 U3724 (.IN1(n7224), .IN2(n2680), .IN3(\key_mem[9][50] ), .IN4(n7212), .Q(n4590)
          );
   AO22X1 U3725 (.IN1(n6804), .IN2(n2680), .IN3(\key_mem[10][50] ), .IN4(n6773), .Q(n4591)
          );
   AO22X1 U3726 (.IN1(n7200), .IN2(n2680), .IN3(\key_mem[11][50] ), .IN4(n7188), .Q(n4592)
          );
   AO22X1 U3727 (.IN1(n7183), .IN2(n2680), .IN3(\key_mem[12][50] ), .IN4(n7184), .Q(n4593)
          );
   AO22X1 U3728 (.IN1(n7179), .IN2(n2680), .IN3(\key_mem[13][50] ), .IN4(n7167), .Q(n4594)
          );
   AO22X1 U3729 (.IN1(n6971), .IN2(n2680), .IN3(\key_mem[14][50] ), .IN4(n7152), .Q(n4595)
          );
   AO222X1 U3731 (.IN1(n7112), .IN2(n2683), .IN3(key[50]), .IN4(n7077), .IN5(n7044), .IN6(
          n2684), .Q(n2682));
   AO22X1 U3732 (.IN1(n7300), .IN2(n2685), .IN3(\key_mem[0][49] ), .IN4(n6932), .Q(n4596)
          );
   AO22X1 U3733 (.IN1(n6810), .IN2(n2685), .IN3(\key_mem[1][49] ), .IN4(n6816), .Q(n4597)
          );
   AO22X1 U3734 (.IN1(n6858), .IN2(n2685), .IN3(\key_mem[2][49] ), .IN4(n6845), .Q(n4598)
          );
   AO22X1 U3735 (.IN1(n6989), .IN2(n2685), .IN3(\key_mem[3][49] ), .IN4(n6864), .Q(n4599)
          );
   AO22X1 U3736 (.IN1(n6990), .IN2(n2685), .IN3(\key_mem[4][49] ), .IN4(n6919), .Q(n4600)
          );
   AO22X1 U3737 (.IN1(n7275), .IN2(n2685), .IN3(\key_mem[5][49] ), .IN4(n7268), .Q(n4601)
          );
   AO22X1 U3738 (.IN1(n7264), .IN2(n2685), .IN3(\key_mem[6][49] ), .IN4(n7015), .Q(n4602)
          );
   AO22X1 U3739 (.IN1(n7250), .IN2(n2685), .IN3(\key_mem[7][49] ), .IN4(n7240), .Q(n4603)
          );
   AO22X1 U3740 (.IN1(n6758), .IN2(n2685), .IN3(\key_mem[8][49] ), .IN4(n6717), .Q(n4604)
          );
   AO22X1 U3741 (.IN1(n7219), .IN2(n2685), .IN3(\key_mem[9][49] ), .IN4(n7213), .Q(n4605)
          );
   AO22X1 U3742 (.IN1(n6805), .IN2(n2685), .IN3(\key_mem[10][49] ), .IN4(n6764), .Q(n4606)
          );
   AO22X1 U3743 (.IN1(n7195), .IN2(n2685), .IN3(\key_mem[11][49] ), .IN4(n7189), .Q(n4607)
          );
   AO22X1 U3744 (.IN1(n6826), .IN2(n2685), .IN3(\key_mem[12][49] ), .IN4(n6985), .Q(n4608)
          );
   AO22X1 U3745 (.IN1(n7174), .IN2(n2685), .IN3(\key_mem[13][49] ), .IN4(n7168), .Q(n4609)
          );
   AO22X1 U3746 (.IN1(n6992), .IN2(n2685), .IN3(\key_mem[14][49] ), .IN4(n7153), .Q(n4610)
          );
   AO221X1 U3747 (.IN1(n7132), .IN2(n2686), .IN3(key[177]), .IN4(n7291), .IN5(n2687), .Q(
          n2685));
   AO222X1 U3748 (.IN1(n7112), .IN2(n2688), .IN3(key[49]), .IN4(n7077), .IN5(n7044), .IN6(
          n2689), .Q(n2687));
   AO22X1 U3749 (.IN1(n7308), .IN2(n2690), .IN3(\key_mem[0][48] ), .IN4(n6932), .Q(n4611)
          );
   AO22X1 U3750 (.IN1(n6813), .IN2(n2690), .IN3(\key_mem[1][48] ), .IN4(n6816), .Q(n4612)
          );
   AO22X1 U3751 (.IN1(n6853), .IN2(n2690), .IN3(\key_mem[2][48] ), .IN4(n6843), .Q(n4613)
          );
   AO22X1 U3752 (.IN1(n6872), .IN2(n2690), .IN3(\key_mem[3][48] ), .IN4(n6876), .Q(n4614)
          );
   AO22X1 U3753 (.IN1(n6916), .IN2(n2690), .IN3(\key_mem[4][48] ), .IN4(n6918), .Q(n4615)
          );
   AO22X1 U3754 (.IN1(n6973), .IN2(n2690), .IN3(\key_mem[5][48] ), .IN4(n7281), .Q(n4616)
          );
   AO22X1 U3755 (.IN1(n7263), .IN2(n2690), .IN3(\key_mem[6][48] ), .IN4(n7253), .Q(n4617)
          );
   AO22X1 U3756 (.IN1(n7249), .IN2(n2690), .IN3(\key_mem[7][48] ), .IN4(n2284), .Q(n4618)
          );
   AO22X1 U3757 (.IN1(n6748), .IN2(n2690), .IN3(\key_mem[8][48] ), .IN4(n6717), .Q(n4619)
          );
   AO22X1 U3758 (.IN1(n6975), .IN2(n2690), .IN3(\key_mem[9][48] ), .IN4(n7225), .Q(n4620)
          );
   AO22X1 U3759 (.IN1(n6795), .IN2(n2690), .IN3(\key_mem[10][48] ), .IN4(n6764), .Q(n4621)
          );
   AO22X1 U3760 (.IN1(n6977), .IN2(n2690), .IN3(\key_mem[11][48] ), .IN4(n7201), .Q(n4622)
          );
   AO22X1 U3761 (.IN1(n7183), .IN2(n2690), .IN3(\key_mem[12][48] ), .IN4(n6828), .Q(n4623)
          );
   AO22X1 U3762 (.IN1(n6979), .IN2(n2690), .IN3(\key_mem[13][48] ), .IN4(n7180), .Q(n4624)
          );
   AO22X1 U3763 (.IN1(n6971), .IN2(n2690), .IN3(\key_mem[14][48] ), .IN4(n7150), .Q(n4625)
          );
   AO221X1 U3764 (.IN1(n7132), .IN2(n2691), .IN3(key[176]), .IN4(n7290), .IN5(n2692), .Q(
          n2690));
   AO222X1 U3765 (.IN1(n7112), .IN2(n2693), .IN3(key[48]), .IN4(n7077), .IN5(n7044), .IN6(
          n2694), .Q(n2692));
   AO22X1 U3766 (.IN1(n7307), .IN2(n2695), .IN3(\key_mem[0][47] ), .IN4(n6931), .Q(n4626)
          );
   AO22X1 U3767 (.IN1(n6810), .IN2(n2695), .IN3(\key_mem[1][47] ), .IN4(n6817), .Q(n4627)
          );
   AO22X1 U3768 (.IN1(n6988), .IN2(n2695), .IN3(\key_mem[2][47] ), .IN4(n6848), .Q(n4628)
          );
   AO22X1 U3769 (.IN1(n6871), .IN2(n2695), .IN3(\key_mem[3][47] ), .IN4(n6863), .Q(n4629)
          );
   AO22X1 U3770 (.IN1(n6924), .IN2(n2695), .IN3(\key_mem[4][47] ), .IN4(n6918), .Q(n4630)
          );
   AO22X1 U3771 (.IN1(n7279), .IN2(n2695), .IN3(\key_mem[5][47] ), .IN4(n7018), .Q(n4631)
          );
   AO22X1 U3772 (.IN1(n7262), .IN2(n2695), .IN3(\key_mem[6][47] ), .IN4(n7251), .Q(n4632)
          );
   AO22X1 U3773 (.IN1(n7013), .IN2(n2695), .IN3(\key_mem[7][47] ), .IN4(n7241), .Q(n4633)
          );
   AO22X1 U3774 (.IN1(n6749), .IN2(n2695), .IN3(\key_mem[8][47] ), .IN4(n6733), .Q(n4634)
          );
   AO22X1 U3775 (.IN1(n7223), .IN2(n2695), .IN3(\key_mem[9][47] ), .IN4(n7007), .Q(n4635)
          );
   AO22X1 U3776 (.IN1(n6796), .IN2(n2695), .IN3(\key_mem[10][47] ), .IN4(n6780), .Q(n4636)
          );
   AO22X1 U3777 (.IN1(n7199), .IN2(n2695), .IN3(\key_mem[11][47] ), .IN4(n7002), .Q(n4637)
          );
   AO22X1 U3778 (.IN1(n6840), .IN2(n2695), .IN3(\key_mem[12][47] ), .IN4(n6983), .Q(n4638)
          );
   AO22X1 U3779 (.IN1(n7178), .IN2(n2695), .IN3(\key_mem[13][47] ), .IN4(n6997), .Q(n4639)
          );
   AO22X1 U3780 (.IN1(n7163), .IN2(n2695), .IN3(\key_mem[14][47] ), .IN4(n7151), .Q(n4640)
          );
   AO221X1 U3781 (.IN1(n7132), .IN2(n2696), .IN3(key[175]), .IN4(n7291), .IN5(n2697), .Q(
          n2695));
   AO222X1 U3782 (.IN1(n7112), .IN2(n2698), .IN3(key[47]), .IN4(n7077), .IN5(n7044), .IN6(
          n2699), .Q(n2697));
   AO22X1 U3783 (.IN1(n7306), .IN2(n2700), .IN3(\key_mem[0][46] ), .IN4(n6931), .Q(n4641)
          );
   AO22X1 U3784 (.IN1(n6927), .IN2(n2700), .IN3(\key_mem[1][46] ), .IN4(n6822), .Q(n4642)
          );
   AO22X1 U3785 (.IN1(n6852), .IN2(n2700), .IN3(\key_mem[2][46] ), .IN4(n6847), .Q(n4643)
          );
   AO22X1 U3786 (.IN1(n6872), .IN2(n2700), .IN3(\key_mem[3][46] ), .IN4(n6864), .Q(n4644)
          );
   AO22X1 U3787 (.IN1(n6920), .IN2(n2700), .IN3(\key_mem[4][46] ), .IN4(n6918), .Q(n4645)
          );
   AO22X1 U3788 (.IN1(n6973), .IN2(n2700), .IN3(\key_mem[5][46] ), .IN4(n7268), .Q(n4646)
          );
   AO22X1 U3789 (.IN1(n7266), .IN2(n2700), .IN3(\key_mem[6][46] ), .IN4(n7251), .Q(n4647)
          );
   AO22X1 U3790 (.IN1(n7250), .IN2(n2700), .IN3(\key_mem[7][46] ), .IN4(n7237), .Q(n4648)
          );
   AO22X1 U3791 (.IN1(n6750), .IN2(n2700), .IN3(\key_mem[8][46] ), .IN4(n6734), .Q(n4649)
          );
   AO22X1 U3792 (.IN1(n6975), .IN2(n2700), .IN3(\key_mem[9][46] ), .IN4(n7212), .Q(n4650)
          );
   AO22X1 U3793 (.IN1(n6797), .IN2(n2700), .IN3(\key_mem[10][46] ), .IN4(n6781), .Q(n4651)
          );
   AO22X1 U3794 (.IN1(n6977), .IN2(n2700), .IN3(\key_mem[11][46] ), .IN4(n7188), .Q(n4652)
          );
   AO22X1 U3795 (.IN1(n6827), .IN2(n2700), .IN3(\key_mem[12][46] ), .IN4(n6833), .Q(n4653)
          );
   AO22X1 U3796 (.IN1(n6979), .IN2(n2700), .IN3(\key_mem[13][46] ), .IN4(n7167), .Q(n4654)
          );
   AO22X1 U3797 (.IN1(n7159), .IN2(n2700), .IN3(\key_mem[14][46] ), .IN4(n7152), .Q(n4655)
          );
   AO221X1 U3798 (.IN1(n7132), .IN2(n2701), .IN3(key[174]), .IN4(n7296), .IN5(n2702), .Q(
          n2700));
   AO222X1 U3799 (.IN1(n7112), .IN2(n2703), .IN3(key[46]), .IN4(n7077), .IN5(n7044), .IN6(
          n2704), .Q(n2702));
   AO22X1 U3800 (.IN1(n7305), .IN2(n2705), .IN3(\key_mem[0][45] ), .IN4(n6931), .Q(n4656)
          );
   AO22X1 U3801 (.IN1(n6812), .IN2(n2705), .IN3(\key_mem[1][45] ), .IN4(n6825), .Q(n4657)
          );
   AO22X1 U3802 (.IN1(n6857), .IN2(n2705), .IN3(\key_mem[2][45] ), .IN4(n6849), .Q(n4658)
          );
   AO22X1 U3803 (.IN1(n6871), .IN2(n2705), .IN3(\key_mem[3][45] ), .IN4(n6861), .Q(n4659)
          );
   AO22X1 U3804 (.IN1(n7288), .IN2(n2705), .IN3(\key_mem[4][45] ), .IN4(n6914), .Q(n4660)
          );
   AO22X1 U3805 (.IN1(n7019), .IN2(n2705), .IN3(\key_mem[5][45] ), .IN4(n7268), .Q(n4661)
          );
   AO22X1 U3806 (.IN1(n7260), .IN2(n2705), .IN3(\key_mem[6][45] ), .IN4(n7251), .Q(n4662)
          );
   AO22X1 U3807 (.IN1(n7250), .IN2(n2705), .IN3(\key_mem[7][45] ), .IN4(n7235), .Q(n4663)
          );
   AO22X1 U3808 (.IN1(n6757), .IN2(n2705), .IN3(\key_mem[8][45] ), .IN4(n6721), .Q(n4664)
          );
   AO22X1 U3809 (.IN1(n7008), .IN2(n2705), .IN3(\key_mem[9][45] ), .IN4(n7213), .Q(n4665)
          );
   AO22X1 U3810 (.IN1(n6804), .IN2(n2705), .IN3(\key_mem[10][45] ), .IN4(n6768), .Q(n4666)
          );
   AO22X1 U3811 (.IN1(n7003), .IN2(n2705), .IN3(\key_mem[11][45] ), .IN4(n7189), .Q(n4667)
          );
   AO22X1 U3812 (.IN1(n6826), .IN2(n2705), .IN3(\key_mem[12][45] ), .IN4(n6839), .Q(n4668)
          );
   AO22X1 U3813 (.IN1(n6998), .IN2(n2705), .IN3(\key_mem[13][45] ), .IN4(n7168), .Q(n4669)
          );
   AO22X1 U3814 (.IN1(n7163), .IN2(n2705), .IN3(\key_mem[14][45] ), .IN4(n7153), .Q(n4670)
          );
   AO221X1 U3815 (.IN1(n7132), .IN2(n2706), .IN3(key[173]), .IN4(n7291), .IN5(n2707), .Q(
          n2705));
   AO222X1 U3816 (.IN1(n7112), .IN2(n2708), .IN3(key[45]), .IN4(n7077), .IN5(n7044), .IN6(
          n2709), .Q(n2707));
   AO22X1 U3817 (.IN1(n7309), .IN2(n2710), .IN3(\key_mem[0][44] ), .IN4(n6931), .Q(n4671)
          );
   AO22X1 U3818 (.IN1(n6810), .IN2(n2710), .IN3(\key_mem[1][44] ), .IN4(n6823), .Q(n4672)
          );
   AO22X1 U3819 (.IN1(n6857), .IN2(n2710), .IN3(\key_mem[2][44] ), .IN4(n6859), .Q(n4673)
          );
   AO22X1 U3820 (.IN1(n6989), .IN2(n2710), .IN3(\key_mem[3][44] ), .IN4(n6868), .Q(n4674)
          );
   AO22X1 U3821 (.IN1(n6924), .IN2(n2710), .IN3(\key_mem[4][44] ), .IN4(n6914), .Q(n4675)
          );
   AO22X1 U3822 (.IN1(n7278), .IN2(n2710), .IN3(\key_mem[5][44] ), .IN4(n7267), .Q(n4676)
          );
   AO22X1 U3823 (.IN1(n7265), .IN2(n2710), .IN3(\key_mem[6][44] ), .IN4(n7259), .Q(n4677)
          );
   AO22X1 U3824 (.IN1(n7246), .IN2(n2710), .IN3(\key_mem[7][44] ), .IN4(n7238), .Q(n4678)
          );
   AO22X1 U3825 (.IN1(n6758), .IN2(n2710), .IN3(\key_mem[8][44] ), .IN4(n7228), .Q(n4679)
          );
   AO22X1 U3826 (.IN1(n7222), .IN2(n2710), .IN3(\key_mem[9][44] ), .IN4(n7211), .Q(n4680)
          );
   AO22X1 U3827 (.IN1(n6805), .IN2(n2710), .IN3(\key_mem[10][44] ), .IN4(n7204), .Q(n4681)
          );
   AO22X1 U3828 (.IN1(n7198), .IN2(n2710), .IN3(\key_mem[11][44] ), .IN4(n7187), .Q(n4682)
          );
   AO22X1 U3829 (.IN1(n6987), .IN2(n2710), .IN3(\key_mem[12][44] ), .IN4(n6833), .Q(n4683)
          );
   AO22X1 U3830 (.IN1(n7177), .IN2(n2710), .IN3(\key_mem[13][44] ), .IN4(n7166), .Q(n4684)
          );
   AO22X1 U3831 (.IN1(n6972), .IN2(n2710), .IN3(\key_mem[14][44] ), .IN4(n7150), .Q(n4685)
          );
   AO221X1 U3832 (.IN1(n7132), .IN2(n2711), .IN3(key[172]), .IN4(n7309), .IN5(n2712), .Q(
          n2710));
   AO222X1 U3833 (.IN1(n7112), .IN2(n2713), .IN3(key[44]), .IN4(n7077), .IN5(n7044), .IN6(
          n2714), .Q(n2712));
   AO22X1 U3834 (.IN1(n7307), .IN2(n2715), .IN3(\key_mem[0][43] ), .IN4(n6931), .Q(n4686)
          );
   AO22X1 U3835 (.IN1(n6812), .IN2(n2715), .IN3(\key_mem[1][43] ), .IN4(n6824), .Q(n4687)
          );
   AO22X1 U3836 (.IN1(n6857), .IN2(n2715), .IN3(\key_mem[2][43] ), .IN4(n6842), .Q(n4688)
          );
   AO22X1 U3837 (.IN1(n6873), .IN2(n2715), .IN3(\key_mem[3][43] ), .IN4(n6867), .Q(n4689)
          );
   AO22X1 U3838 (.IN1(n6889), .IN2(n2715), .IN3(\key_mem[4][43] ), .IN4(n6915), .Q(n4690)
          );
   AO22X1 U3839 (.IN1(n7019), .IN2(n2715), .IN3(\key_mem[5][43] ), .IN4(n7267), .Q(n4691)
          );
   AO22X1 U3840 (.IN1(n7260), .IN2(n2715), .IN3(\key_mem[6][43] ), .IN4(n7257), .Q(n4692)
          );
   AO22X1 U3841 (.IN1(n7249), .IN2(n2715), .IN3(\key_mem[7][43] ), .IN4(n7012), .Q(n4693)
          );
   AO22X1 U3842 (.IN1(n6748), .IN2(n2715), .IN3(\key_mem[8][43] ), .IN4(n6721), .Q(n4694)
          );
   AO22X1 U3843 (.IN1(n7008), .IN2(n2715), .IN3(\key_mem[9][43] ), .IN4(n7211), .Q(n4695)
          );
   AO22X1 U3844 (.IN1(n6795), .IN2(n2715), .IN3(\key_mem[10][43] ), .IN4(n6768), .Q(n4696)
          );
   AO22X1 U3845 (.IN1(n7003), .IN2(n2715), .IN3(\key_mem[11][43] ), .IN4(n7187), .Q(n4697)
          );
   AO22X1 U3846 (.IN1(n7001), .IN2(n2715), .IN3(\key_mem[12][43] ), .IN4(n6982), .Q(n4698)
          );
   AO22X1 U3847 (.IN1(n6998), .IN2(n2715), .IN3(\key_mem[13][43] ), .IN4(n7166), .Q(n4699)
          );
   AO22X1 U3848 (.IN1(n7163), .IN2(n2715), .IN3(\key_mem[14][43] ), .IN4(n7151), .Q(n4700)
          );
   AO221X1 U3849 (.IN1(n7133), .IN2(n2716), .IN3(key[171]), .IN4(n7312), .IN5(n2717), .Q(
          n2715));
   AO222X1 U3850 (.IN1(n7111), .IN2(n2718), .IN3(key[43]), .IN4(n7078), .IN5(n7045), .IN6(
          n2719), .Q(n2717));
   AO22X1 U3851 (.IN1(n7304), .IN2(n2720), .IN3(\key_mem[0][42] ), .IN4(n6931), .Q(n4701)
          );
   AO22X1 U3852 (.IN1(n6926), .IN2(n2720), .IN3(\key_mem[1][42] ), .IN4(n6825), .Q(n4702)
          );
   AO22X1 U3853 (.IN1(n6854), .IN2(n2720), .IN3(\key_mem[2][42] ), .IN4(n6850), .Q(n4703)
          );
   AO22X1 U3854 (.IN1(n6989), .IN2(n2720), .IN3(\key_mem[3][42] ), .IN4(n6862), .Q(n4704)
          );
   AO22X1 U3855 (.IN1(n7287), .IN2(n2720), .IN3(\key_mem[4][42] ), .IN4(n6917), .Q(n4705)
          );
   AO22X1 U3856 (.IN1(n7020), .IN2(n2720), .IN3(\key_mem[5][42] ), .IN4(n7281), .Q(n4706)
          );
   AO22X1 U3857 (.IN1(n7260), .IN2(n2720), .IN3(\key_mem[6][42] ), .IN4(n7251), .Q(n4707)
          );
   AO22X1 U3858 (.IN1(n7014), .IN2(n2720), .IN3(\key_mem[7][42] ), .IN4(n7243), .Q(n4708)
          );
   AO22X1 U3859 (.IN1(n6749), .IN2(n2720), .IN3(\key_mem[8][42] ), .IN4(n6719), .Q(n4709)
          );
   AO22X1 U3860 (.IN1(n7009), .IN2(n2720), .IN3(\key_mem[9][42] ), .IN4(n7225), .Q(n4710)
          );
   AO22X1 U3861 (.IN1(n6796), .IN2(n2720), .IN3(\key_mem[10][42] ), .IN4(n6766), .Q(n4711)
          );
   AO22X1 U3862 (.IN1(n7004), .IN2(n2720), .IN3(\key_mem[11][42] ), .IN4(n7201), .Q(n4712)
          );
   AO22X1 U3863 (.IN1(n7186), .IN2(n2720), .IN3(\key_mem[12][42] ), .IN4(n7185), .Q(n4713)
          );
   AO22X1 U3864 (.IN1(n6999), .IN2(n2720), .IN3(\key_mem[13][42] ), .IN4(n7180), .Q(n4714)
          );
   AO22X1 U3865 (.IN1(n6972), .IN2(n2720), .IN3(\key_mem[14][42] ), .IN4(n7150), .Q(n4715)
          );
   AO222X1 U3867 (.IN1(n7111), .IN2(n2723), .IN3(key[42]), .IN4(n7078), .IN5(n7045), .IN6(
          n2724), .Q(n2722));
   AO22X1 U3868 (.IN1(n7312), .IN2(n2725), .IN3(\key_mem[0][41] ), .IN4(n6931), .Q(n4716)
          );
   AO22X1 U3869 (.IN1(n6926), .IN2(n2725), .IN3(\key_mem[1][41] ), .IN4(n6820), .Q(n4717)
          );
   AO22X1 U3870 (.IN1(n6855), .IN2(n2725), .IN3(\key_mem[2][41] ), .IN4(n6844), .Q(n4718)
          );
   AO22X1 U3871 (.IN1(n6872), .IN2(n2725), .IN3(\key_mem[3][41] ), .IN4(n6877), .Q(n4719)
          );
   AO22X1 U3872 (.IN1(n6920), .IN2(n2725), .IN3(\key_mem[4][41] ), .IN4(n6923), .Q(n4720)
          );
   AO22X1 U3873 (.IN1(n7278), .IN2(n2725), .IN3(\key_mem[5][41] ), .IN4(n7282), .Q(n4721)
          );
   AO22X1 U3874 (.IN1(n7260), .IN2(n2725), .IN3(\key_mem[6][41] ), .IN4(n7259), .Q(n4722)
          );
   AO22X1 U3875 (.IN1(n7244), .IN2(n2725), .IN3(\key_mem[7][41] ), .IN4(n7235), .Q(n4723)
          );
   AO22X1 U3876 (.IN1(n6750), .IN2(n2725), .IN3(\key_mem[8][41] ), .IN4(n6720), .Q(n4724)
          );
   AO22X1 U3877 (.IN1(n7222), .IN2(n2725), .IN3(\key_mem[9][41] ), .IN4(n7226), .Q(n4725)
          );
   AO22X1 U3878 (.IN1(n6797), .IN2(n2725), .IN3(\key_mem[10][41] ), .IN4(n6767), .Q(n4726)
          );
   AO22X1 U3879 (.IN1(n7198), .IN2(n2725), .IN3(\key_mem[11][41] ), .IN4(n7202), .Q(n4727)
          );
   AO22X1 U3880 (.IN1(n6835), .IN2(n2725), .IN3(\key_mem[12][41] ), .IN4(n6841), .Q(n4728)
          );
   AO22X1 U3881 (.IN1(n7177), .IN2(n2725), .IN3(\key_mem[13][41] ), .IN4(n7181), .Q(n4729)
          );
   AO22X1 U3882 (.IN1(n6971), .IN2(n2725), .IN3(\key_mem[14][41] ), .IN4(n7156), .Q(n4730)
          );
   AO222X1 U3884 (.IN1(n7111), .IN2(n2728), .IN3(key[41]), .IN4(n7078), .IN5(n7045), .IN6(
          n2729), .Q(n2727));
   AO22X1 U3885 (.IN1(n7308), .IN2(n2730), .IN3(\key_mem[0][40] ), .IN4(n6931), .Q(n4731)
          );
   AO22X1 U3886 (.IN1(n6813), .IN2(n2730), .IN3(\key_mem[1][40] ), .IN4(n6820), .Q(n4732)
          );
   AO22X1 U3887 (.IN1(n6858), .IN2(n2730), .IN3(\key_mem[2][40] ), .IN4(n6850), .Q(n4733)
          );
   AO22X1 U3888 (.IN1(n6871), .IN2(n2730), .IN3(\key_mem[3][40] ), .IN4(n6877), .Q(n4734)
          );
   AO22X1 U3889 (.IN1(n7287), .IN2(n2730), .IN3(\key_mem[4][40] ), .IN4(n6914), .Q(n4735)
          );
   AO22X1 U3890 (.IN1(n7280), .IN2(n2730), .IN3(\key_mem[5][40] ), .IN4(n7270), .Q(n4736)
          );
   AO22X1 U3891 (.IN1(n7264), .IN2(n2730), .IN3(\key_mem[6][40] ), .IN4(n7259), .Q(n4737)
          );
   AO22X1 U3892 (.IN1(n7245), .IN2(n2730), .IN3(\key_mem[7][40] ), .IN4(n7236), .Q(n4738)
          );
   AO22X1 U3893 (.IN1(n6749), .IN2(n2730), .IN3(\key_mem[8][40] ), .IN4(n6720), .Q(n4739)
          );
   AO22X1 U3894 (.IN1(n7224), .IN2(n2730), .IN3(\key_mem[9][40] ), .IN4(n7212), .Q(n4740)
          );
   AO22X1 U3895 (.IN1(n6796), .IN2(n2730), .IN3(\key_mem[10][40] ), .IN4(n6767), .Q(n4741)
          );
   AO22X1 U3896 (.IN1(n7200), .IN2(n2730), .IN3(\key_mem[11][40] ), .IN4(n7188), .Q(n4742)
          );
   AO22X1 U3897 (.IN1(n7001), .IN2(n2730), .IN3(\key_mem[12][40] ), .IN4(n6982), .Q(n4743)
          );
   AO22X1 U3898 (.IN1(n7179), .IN2(n2730), .IN3(\key_mem[13][40] ), .IN4(n7167), .Q(n4744)
          );
   AO22X1 U3899 (.IN1(n6995), .IN2(n2730), .IN3(\key_mem[14][40] ), .IN4(n7147), .Q(n4745)
          );
   AO221X1 U3900 (.IN1(n7133), .IN2(n2731), .IN3(key[168]), .IN4(n7293), .IN5(n2732), .Q(
          n2730));
   AO222X1 U3901 (.IN1(n7111), .IN2(n2733), .IN3(key[40]), .IN4(n7078), .IN5(n7045), .IN6(
          n2734), .Q(n2732));
   AO22X1 U3902 (.IN1(n7307), .IN2(n2735), .IN3(\key_mem[0][39] ), .IN4(n6931), .Q(n4746)
          );
   AO22X1 U3903 (.IN1(n6808), .IN2(n2735), .IN3(\key_mem[1][39] ), .IN4(n6818), .Q(n4747)
          );
   AO22X1 U3904 (.IN1(n6853), .IN2(n2735), .IN3(\key_mem[2][39] ), .IN4(n6849), .Q(n4748)
          );
   AO22X1 U3905 (.IN1(n6807), .IN2(n2735), .IN3(\key_mem[3][39] ), .IN4(n6861), .Q(n4749)
          );
   AO22X1 U3906 (.IN1(n6888), .IN2(n2735), .IN3(\key_mem[4][39] ), .IN4(n6923), .Q(n4750)
          );
   AO22X1 U3907 (.IN1(n7279), .IN2(n2735), .IN3(\key_mem[5][39] ), .IN4(n7267), .Q(n4751)
          );
   AO22X1 U3908 (.IN1(n7261), .IN2(n2735), .IN3(\key_mem[6][39] ), .IN4(n7258), .Q(n4752)
          );
   AO22X1 U3909 (.IN1(n7246), .IN2(n2735), .IN3(\key_mem[7][39] ), .IN4(n7237), .Q(n4753)
          );
   AO22X1 U3910 (.IN1(n6750), .IN2(n2735), .IN3(\key_mem[8][39] ), .IN4(n6718), .Q(n4754)
          );
   AO22X1 U3911 (.IN1(n7223), .IN2(n2735), .IN3(\key_mem[9][39] ), .IN4(n7211), .Q(n4755)
          );
   AO22X1 U3912 (.IN1(n6797), .IN2(n2735), .IN3(\key_mem[10][39] ), .IN4(n6765), .Q(n4756)
          );
   AO22X1 U3913 (.IN1(n7199), .IN2(n2735), .IN3(\key_mem[11][39] ), .IN4(n7187), .Q(n4757)
          );
   AO22X1 U3914 (.IN1(n6831), .IN2(n2735), .IN3(\key_mem[12][39] ), .IN4(n7185), .Q(n4758)
          );
   AO22X1 U3915 (.IN1(n7178), .IN2(n2735), .IN3(\key_mem[13][39] ), .IN4(n7166), .Q(n4759)
          );
   AO22X1 U3916 (.IN1(n7164), .IN2(n2735), .IN3(\key_mem[14][39] ), .IN4(n7153), .Q(n4760)
          );
   AO221X1 U3917 (.IN1(n7133), .IN2(n2736), .IN3(key[167]), .IN4(n7291), .IN5(n2737), .Q(
          n2735));
   AO222X1 U3918 (.IN1(n7111), .IN2(n2738), .IN3(key[39]), .IN4(n7078), .IN5(n7045), .IN6(
          n2739), .Q(n2737));
   AO22X1 U3919 (.IN1(n7306), .IN2(n2740), .IN3(\key_mem[0][38] ), .IN4(n6931), .Q(n4761)
          );
   AO22X1 U3920 (.IN1(n6813), .IN2(n2740), .IN3(\key_mem[1][38] ), .IN4(n6819), .Q(n4762)
          );
   AO22X1 U3921 (.IN1(n6858), .IN2(n2740), .IN3(\key_mem[2][38] ), .IN4(n6844), .Q(n4763)
          );
   AO22X1 U3922 (.IN1(n6989), .IN2(n2740), .IN3(\key_mem[3][38] ), .IN4(n6877), .Q(n4764)
          );
   AO22X1 U3923 (.IN1(n6886), .IN2(n2740), .IN3(\key_mem[4][38] ), .IN4(n6919), .Q(n4765)
          );
   AO22X1 U3924 (.IN1(n7274), .IN2(n2740), .IN3(\key_mem[5][38] ), .IN4(n7269), .Q(n4766)
          );
   AO22X1 U3925 (.IN1(n7260), .IN2(n2740), .IN3(\key_mem[6][38] ), .IN4(n7256), .Q(n4767)
          );
   AO22X1 U3926 (.IN1(n7247), .IN2(n2740), .IN3(\key_mem[7][38] ), .IN4(n7238), .Q(n4768)
          );
   AO22X1 U3927 (.IN1(n6751), .IN2(n2740), .IN3(\key_mem[8][38] ), .IN4(n6714), .Q(n4769)
          );
   AO22X1 U3928 (.IN1(n7218), .IN2(n2740), .IN3(\key_mem[9][38] ), .IN4(n7212), .Q(n4770)
          );
   AO22X1 U3929 (.IN1(n6798), .IN2(n2740), .IN3(\key_mem[10][38] ), .IN4(n6761), .Q(n4771)
          );
   AO22X1 U3930 (.IN1(n7194), .IN2(n2740), .IN3(\key_mem[11][38] ), .IN4(n7188), .Q(n4772)
          );
   AO22X1 U3931 (.IN1(n7183), .IN2(n2740), .IN3(\key_mem[12][38] ), .IN4(n7000), .Q(n4773)
          );
   AO22X1 U3932 (.IN1(n7173), .IN2(n2740), .IN3(\key_mem[13][38] ), .IN4(n7167), .Q(n4774)
          );
   AO22X1 U3933 (.IN1(n6996), .IN2(n2740), .IN3(\key_mem[14][38] ), .IN4(n7148), .Q(n4775)
          );
   AO222X1 U3935 (.IN1(n7111), .IN2(n2743), .IN3(key[38]), .IN4(n7078), .IN5(n7045), .IN6(
          n2744), .Q(n2742));
   AO22X1 U3936 (.IN1(n7305), .IN2(n2745), .IN3(\key_mem[0][37] ), .IN4(n6931), .Q(n4776)
          );
   AO22X1 U3937 (.IN1(n6812), .IN2(n2745), .IN3(\key_mem[1][37] ), .IN4(n6817), .Q(n4777)
          );
   AO22X1 U3938 (.IN1(n6854), .IN2(n2745), .IN3(\key_mem[2][37] ), .IN4(n6850), .Q(n4778)
          );
   AO22X1 U3939 (.IN1(n6874), .IN2(n2745), .IN3(\key_mem[3][37] ), .IN4(n6866), .Q(n4779)
          );
   AO22X1 U3940 (.IN1(n6887), .IN2(n2745), .IN3(\key_mem[4][37] ), .IN4(n6918), .Q(n4780)
          );
   AO22X1 U3941 (.IN1(n7276), .IN2(n2745), .IN3(\key_mem[5][37] ), .IN4(n7269), .Q(n4781)
          );
   AO22X1 U3942 (.IN1(n7265), .IN2(n2745), .IN3(\key_mem[6][37] ), .IN4(n7257), .Q(n4782)
          );
   AO22X1 U3943 (.IN1(n7249), .IN2(n2745), .IN3(\key_mem[7][37] ), .IN4(n7239), .Q(n4783)
          );
   AO22X1 U3944 (.IN1(n6751), .IN2(n2745), .IN3(\key_mem[8][37] ), .IN4(n6715), .Q(n4784)
          );
   AO22X1 U3945 (.IN1(n7220), .IN2(n2745), .IN3(\key_mem[9][37] ), .IN4(n7214), .Q(n4785)
          );
   AO22X1 U3946 (.IN1(n6798), .IN2(n2745), .IN3(\key_mem[10][37] ), .IN4(n6762), .Q(n4786)
          );
   AO22X1 U3947 (.IN1(n7196), .IN2(n2745), .IN3(\key_mem[11][37] ), .IN4(n7190), .Q(n4787)
          );
   AO22X1 U3948 (.IN1(n6826), .IN2(n2745), .IN3(\key_mem[12][37] ), .IN4(n6983), .Q(n4788)
          );
   AO22X1 U3949 (.IN1(n7175), .IN2(n2745), .IN3(\key_mem[13][37] ), .IN4(n7169), .Q(n4789)
          );
   AO22X1 U3950 (.IN1(n7159), .IN2(n2745), .IN3(\key_mem[14][37] ), .IN4(n7149), .Q(n4790)
          );
   AO221X1 U3951 (.IN1(n7133), .IN2(n2746), .IN3(key[165]), .IN4(n7293), .IN5(n2747), .Q(
          n2745));
   AO222X1 U3952 (.IN1(n7111), .IN2(n2748), .IN3(key[37]), .IN4(n7078), .IN5(n7045), .IN6(
          n2749), .Q(n2747));
   AO22X1 U3953 (.IN1(n7309), .IN2(n2750), .IN3(\key_mem[0][36] ), .IN4(n6931), .Q(n4791)
          );
   AO22X1 U3954 (.IN1(n6809), .IN2(n2750), .IN3(\key_mem[1][36] ), .IN4(n6818), .Q(n4792)
          );
   AO22X1 U3955 (.IN1(n6854), .IN2(n2750), .IN3(\key_mem[2][36] ), .IN4(n6842), .Q(n4793)
          );
   AO22X1 U3956 (.IN1(n6874), .IN2(n2750), .IN3(\key_mem[3][36] ), .IN4(n6876), .Q(n4794)
          );
   AO22X1 U3957 (.IN1(n7286), .IN2(n2750), .IN3(\key_mem[4][36] ), .IN4(n7285), .Q(n4795)
          );
   AO22X1 U3958 (.IN1(n7283), .IN2(n2750), .IN3(\key_mem[5][36] ), .IN4(n7270), .Q(n4796)
          );
   AO22X1 U3959 (.IN1(n6970), .IN2(n2750), .IN3(\key_mem[6][36] ), .IN4(n7254), .Q(n4797)
          );
   AO22X1 U3960 (.IN1(n7249), .IN2(n2750), .IN3(\key_mem[7][36] ), .IN4(n7240), .Q(n4798)
          );
   AO22X1 U3961 (.IN1(n6752), .IN2(n2750), .IN3(\key_mem[8][36] ), .IN4(n6716), .Q(n4799)
          );
   AO22X1 U3962 (.IN1(n7227), .IN2(n2750), .IN3(\key_mem[9][36] ), .IN4(n7214), .Q(n4800)
          );
   AO22X1 U3963 (.IN1(n6799), .IN2(n2750), .IN3(\key_mem[10][36] ), .IN4(n6763), .Q(n4801)
          );
   AO22X1 U3964 (.IN1(n7203), .IN2(n2750), .IN3(\key_mem[11][36] ), .IN4(n7190), .Q(n4802)
          );
   AO22X1 U3965 (.IN1(n6986), .IN2(n2750), .IN3(\key_mem[12][36] ), .IN4(n6984), .Q(n4803)
          );
   AO22X1 U3966 (.IN1(n7182), .IN2(n2750), .IN3(\key_mem[13][36] ), .IN4(n7169), .Q(n4804)
          );
   AO22X1 U3967 (.IN1(n6992), .IN2(n2750), .IN3(\key_mem[14][36] ), .IN4(n7156), .Q(n4805)
          );
   AO221X1 U3968 (.IN1(n7133), .IN2(n2751), .IN3(key[164]), .IN4(n7290), .IN5(n2752), .Q(
          n2750));
   AO222X1 U3969 (.IN1(n7111), .IN2(n2753), .IN3(key[36]), .IN4(n7078), .IN5(n7045), .IN6(
          n2754), .Q(n2752));
   AO22X1 U3970 (.IN1(n7311), .IN2(n2755), .IN3(\key_mem[0][35] ), .IN4(n6930), .Q(n4806)
          );
   AO22X1 U3971 (.IN1(n6809), .IN2(n2755), .IN3(\key_mem[1][35] ), .IN4(n6822), .Q(n4807)
          );
   AO22X1 U3972 (.IN1(n6856), .IN2(n2755), .IN3(\key_mem[2][35] ), .IN4(n6851), .Q(n4808)
          );
   AO22X1 U3973 (.IN1(n6875), .IN2(n2755), .IN3(\key_mem[3][35] ), .IN4(n6877), .Q(n4809)
          );
   AO22X1 U3974 (.IN1(n6924), .IN2(n2755), .IN3(\key_mem[4][35] ), .IN4(n6917), .Q(n4810)
          );
   AO22X1 U3975 (.IN1(n6974), .IN2(n2755), .IN3(\key_mem[5][35] ), .IN4(n7268), .Q(n4811)
          );
   AO22X1 U3976 (.IN1(n7264), .IN2(n2755), .IN3(\key_mem[6][35] ), .IN4(n7015), .Q(n4812)
          );
   AO22X1 U3977 (.IN1(n7247), .IN2(n2755), .IN3(\key_mem[7][35] ), .IN4(n7241), .Q(n4813)
          );
   AO22X1 U3978 (.IN1(n6749), .IN2(n2755), .IN3(\key_mem[8][35] ), .IN4(n6725), .Q(n4814)
          );
   AO22X1 U3979 (.IN1(n6976), .IN2(n2755), .IN3(\key_mem[9][35] ), .IN4(n7213), .Q(n4815)
          );
   AO22X1 U3980 (.IN1(n6796), .IN2(n2755), .IN3(\key_mem[10][35] ), .IN4(n6772), .Q(n4816)
          );
   AO22X1 U3981 (.IN1(n6978), .IN2(n2755), .IN3(\key_mem[11][35] ), .IN4(n7189), .Q(n4817)
          );
   AO22X1 U3982 (.IN1(n6835), .IN2(n2755), .IN3(\key_mem[12][35] ), .IN4(n6838), .Q(n4818)
          );
   AO22X1 U3983 (.IN1(n6980), .IN2(n2755), .IN3(\key_mem[13][35] ), .IN4(n7168), .Q(n4819)
          );
   AO22X1 U3984 (.IN1(n6972), .IN2(n2755), .IN3(\key_mem[14][35] ), .IN4(n7151), .Q(n4820)
          );
   AO221X1 U3985 (.IN1(n7133), .IN2(n2756), .IN3(key[163]), .IN4(n7291), .IN5(n2757), .Q(
          n2755));
   AO222X1 U3986 (.IN1(n7111), .IN2(n2758), .IN3(key[35]), .IN4(n7078), .IN5(n7045), .IN6(
          n2759), .Q(n2757));
   AO22X1 U3987 (.IN1(n7312), .IN2(n2760), .IN3(\key_mem[0][34] ), .IN4(n6930), .Q(n4821)
          );
   AO22X1 U3988 (.IN1(n6811), .IN2(n2760), .IN3(\key_mem[1][34] ), .IN4(n6816), .Q(n4822)
          );
   AO22X1 U3989 (.IN1(n6988), .IN2(n2760), .IN3(\key_mem[2][34] ), .IN4(n6851), .Q(n4823)
          );
   AO22X1 U3990 (.IN1(n6807), .IN2(n2760), .IN3(\key_mem[3][34] ), .IN4(n6860), .Q(n4824)
          );
   AO22X1 U3991 (.IN1(n6924), .IN2(n2760), .IN3(\key_mem[4][34] ), .IN4(n6915), .Q(n4825)
          );
   AO22X1 U3992 (.IN1(n7283), .IN2(n2760), .IN3(\key_mem[5][34] ), .IN4(n7272), .Q(n4826)
          );
   AO22X1 U3993 (.IN1(n6970), .IN2(n2760), .IN3(\key_mem[6][34] ), .IN4(n7259), .Q(n4827)
          );
   AO22X1 U3994 (.IN1(n7013), .IN2(n2760), .IN3(\key_mem[7][34] ), .IN4(n7242), .Q(n4828)
          );
   AO22X1 U3995 (.IN1(n6748), .IN2(n2760), .IN3(\key_mem[8][34] ), .IN4(n6717), .Q(n4829)
          );
   AO22X1 U3996 (.IN1(n7227), .IN2(n2760), .IN3(\key_mem[9][34] ), .IN4(n7215), .Q(n4830)
          );
   AO22X1 U3997 (.IN1(n6795), .IN2(n2760), .IN3(\key_mem[10][34] ), .IN4(n6764), .Q(n4831)
          );
   AO22X1 U3998 (.IN1(n7203), .IN2(n2760), .IN3(\key_mem[11][34] ), .IN4(n7191), .Q(n4832)
          );
   AO22X1 U3999 (.IN1(n6986), .IN2(n2760), .IN3(\key_mem[12][34] ), .IN4(n6836), .Q(n4833)
          );
   AO22X1 U4000 (.IN1(n7182), .IN2(n2760), .IN3(\key_mem[13][34] ), .IN4(n7170), .Q(n4834)
          );
   AO22X1 U4001 (.IN1(n7158), .IN2(n2760), .IN3(\key_mem[14][34] ), .IN4(n7157), .Q(n4835)
          );
   AO221X1 U4002 (.IN1(n7133), .IN2(n2761), .IN3(key[162]), .IN4(n7297), .IN5(n2762), .Q(
          n2760));
   AO222X1 U4003 (.IN1(n7111), .IN2(n2763), .IN3(key[34]), .IN4(n7078), .IN5(n7045), .IN6(
          n2764), .Q(n2762));
   AO22X1 U4004 (.IN1(n2276), .IN2(n2765), .IN3(\key_mem[0][33] ), .IN4(n6930), .Q(n4836)
          );
   AO22X1 U4005 (.IN1(n6811), .IN2(n2765), .IN3(\key_mem[1][33] ), .IN4(n6821), .Q(n4837)
          );
   AO22X1 U4006 (.IN1(n6852), .IN2(n2765), .IN3(\key_mem[2][33] ), .IN4(n6849), .Q(n4838)
          );
   AO22X1 U4007 (.IN1(n6872), .IN2(n2765), .IN3(\key_mem[3][33] ), .IN4(n6867), .Q(n4839)
          );
   AO22X1 U4008 (.IN1(n7288), .IN2(n2765), .IN3(\key_mem[4][33] ), .IN4(n7284), .Q(n4840)
          );
   AO22X1 U4009 (.IN1(n7020), .IN2(n2765), .IN3(\key_mem[5][33] ), .IN4(n7273), .Q(n4841)
          );
   AO22X1 U4010 (.IN1(n6969), .IN2(n2765), .IN3(\key_mem[6][33] ), .IN4(n7252), .Q(n4842)
          );
   AO22X1 U4011 (.IN1(n7248), .IN2(n2765), .IN3(\key_mem[7][33] ), .IN4(n7238), .Q(n4843)
          );
   AO22X1 U4012 (.IN1(n6749), .IN2(n2765), .IN3(\key_mem[8][33] ), .IN4(n6718), .Q(n4844)
          );
   AO22X1 U4013 (.IN1(n7009), .IN2(n2765), .IN3(\key_mem[9][33] ), .IN4(n7217), .Q(n4845)
          );
   AO22X1 U4014 (.IN1(n6796), .IN2(n2765), .IN3(\key_mem[10][33] ), .IN4(n6765), .Q(n4846)
          );
   AO22X1 U4015 (.IN1(n7004), .IN2(n2765), .IN3(\key_mem[11][33] ), .IN4(n7193), .Q(n4847)
          );
   AO22X1 U4016 (.IN1(n6826), .IN2(n2765), .IN3(\key_mem[12][33] ), .IN4(n6838), .Q(n4848)
          );
   AO22X1 U4017 (.IN1(n6999), .IN2(n2765), .IN3(\key_mem[13][33] ), .IN4(n7172), .Q(n4849)
          );
   AO22X1 U4018 (.IN1(n6971), .IN2(n2765), .IN3(\key_mem[14][33] ), .IN4(n6994), .Q(n4850)
          );
   AO222X1 U4020 (.IN1(n7111), .IN2(n2768), .IN3(key[33]), .IN4(n7078), .IN5(n7045), .IN6(
          n2769), .Q(n2767));
   AO22X1 U4021 (.IN1(n7294), .IN2(n2770), .IN3(\key_mem[0][32] ), .IN4(n6930), .Q(n4851)
          );
   AO22X1 U4022 (.IN1(n6809), .IN2(n2770), .IN3(\key_mem[1][32] ), .IN4(n6817), .Q(n4852)
          );
   AO22X1 U4023 (.IN1(n6857), .IN2(n2770), .IN3(\key_mem[2][32] ), .IN4(n6850), .Q(n4853)
          );
   AO22X1 U4024 (.IN1(n6807), .IN2(n2770), .IN3(\key_mem[3][32] ), .IN4(n6863), .Q(n4854)
          );
   AO22X1 U4025 (.IN1(n6889), .IN2(n2770), .IN3(\key_mem[4][32] ), .IN4(n6915), .Q(n4855)
          );
   AO22X1 U4026 (.IN1(n7280), .IN2(n2770), .IN3(\key_mem[5][32] ), .IN4(n7271), .Q(n4856)
          );
   AO22X1 U4027 (.IN1(n7265), .IN2(n2770), .IN3(\key_mem[6][32] ), .IN4(n7253), .Q(n4857)
          );
   AO22X1 U4028 (.IN1(n7250), .IN2(n2770), .IN3(\key_mem[7][32] ), .IN4(n7236), .Q(n4858)
          );
   AO22X1 U4029 (.IN1(n6754), .IN2(n2770), .IN3(\key_mem[8][32] ), .IN4(n6725), .Q(n4859)
          );
   AO22X1 U4030 (.IN1(n7224), .IN2(n2770), .IN3(\key_mem[9][32] ), .IN4(n7215), .Q(n4860)
          );
   AO22X1 U4031 (.IN1(n6801), .IN2(n2770), .IN3(\key_mem[10][32] ), .IN4(n6772), .Q(n4861)
          );
   AO22X1 U4032 (.IN1(n7200), .IN2(n2770), .IN3(\key_mem[11][32] ), .IN4(n7191), .Q(n4862)
          );
   AO22X1 U4033 (.IN1(n7183), .IN2(n2770), .IN3(\key_mem[12][32] ), .IN4(n6838), .Q(n4863)
          );
   AO22X1 U4034 (.IN1(n7179), .IN2(n2770), .IN3(\key_mem[13][32] ), .IN4(n7170), .Q(n4864)
          );
   AO22X1 U4035 (.IN1(n6992), .IN2(n2770), .IN3(\key_mem[14][32] ), .IN4(n7152), .Q(n4865)
          );
   AO221X1 U4036 (.IN1(n7133), .IN2(n2771), .IN3(key[160]), .IN4(n7296), .IN5(n2772), .Q(
          n2770));
   AO222X1 U4037 (.IN1(n7111), .IN2(n2773), .IN3(key[32]), .IN4(n7078), .IN5(n7045), .IN6(
          n2774), .Q(n2772));
   AO22X1 U4038 (.IN1(n7293), .IN2(n2775), .IN3(\key_mem[0][31] ), .IN4(n6930), .Q(n4866)
          );
   AO22X1 U4039 (.IN1(n6808), .IN2(n2775), .IN3(\key_mem[1][31] ), .IN4(n6818), .Q(n4867)
          );
   AO22X1 U4040 (.IN1(n6857), .IN2(n2775), .IN3(\key_mem[2][31] ), .IN4(n6844), .Q(n4868)
          );
   AO22X1 U4041 (.IN1(n6874), .IN2(n2775), .IN3(\key_mem[3][31] ), .IN4(n6876), .Q(n4869)
          );
   AO22X1 U4042 (.IN1(n7287), .IN2(n2775), .IN3(\key_mem[4][31] ), .IN4(n6923), .Q(n4870)
          );
   AO22X1 U4043 (.IN1(n7278), .IN2(n2775), .IN3(\key_mem[5][31] ), .IN4(n7272), .Q(n4871)
          );
   AO22X1 U4044 (.IN1(n7265), .IN2(n2775), .IN3(\key_mem[6][31] ), .IN4(n7255), .Q(n4872)
          );
   AO22X1 U4045 (.IN1(n7249), .IN2(n2775), .IN3(\key_mem[7][31] ), .IN4(n7239), .Q(n4873)
          );
   AO22X1 U4046 (.IN1(n6755), .IN2(n2775), .IN3(\key_mem[8][31] ), .IN4(n6717), .Q(n4874)
          );
   AO22X1 U4047 (.IN1(n7222), .IN2(n2775), .IN3(\key_mem[9][31] ), .IN4(n7216), .Q(n4875)
          );
   AO22X1 U4048 (.IN1(n6802), .IN2(n2775), .IN3(\key_mem[10][31] ), .IN4(n6764), .Q(n4876)
          );
   AO22X1 U4049 (.IN1(n7198), .IN2(n2775), .IN3(\key_mem[11][31] ), .IN4(n7192), .Q(n4877)
          );
   AO22X1 U4050 (.IN1(n6837), .IN2(n2775), .IN3(\key_mem[12][31] ), .IN4(n6982), .Q(n4878)
          );
   AO22X1 U4051 (.IN1(n7177), .IN2(n2775), .IN3(\key_mem[13][31] ), .IN4(n7171), .Q(n4879)
          );
   AO22X1 U4052 (.IN1(n6992), .IN2(n2775), .IN3(\key_mem[14][31] ), .IN4(n7153), .Q(n4880)
          );
   AO221X1 U4053 (.IN1(n7134), .IN2(n2776), .IN3(key[159]), .IN4(n2276), .IN5(n2777), .Q(
          n2775));
   AO222X1 U4054 (.IN1(n7111), .IN2(n2778), .IN3(key[31]), .IN4(n7079), .IN5(n7046), .IN6(
          n2779), .Q(n2777));
   AO22X1 U4055 (.IN1(n7311), .IN2(n2780), .IN3(\key_mem[0][30] ), .IN4(n6930), .Q(n4881)
          );
   AO22X1 U4056 (.IN1(n6812), .IN2(n2780), .IN3(\key_mem[1][30] ), .IN4(n6819), .Q(n4882)
          );
   AO22X1 U4057 (.IN1(n6854), .IN2(n2780), .IN3(\key_mem[2][30] ), .IN4(n6859), .Q(n4883)
          );
   AO22X1 U4058 (.IN1(n6875), .IN2(n2780), .IN3(\key_mem[3][30] ), .IN4(n6867), .Q(n4884)
          );
   AO22X1 U4059 (.IN1(n7288), .IN2(n2780), .IN3(\key_mem[4][30] ), .IN4(n7285), .Q(n4885)
          );
   AO22X1 U4060 (.IN1(n7280), .IN2(n2780), .IN3(\key_mem[5][30] ), .IN4(n7269), .Q(n4886)
          );
   AO22X1 U4061 (.IN1(n7265), .IN2(n2780), .IN3(\key_mem[6][30] ), .IN4(n7252), .Q(n4887)
          );
   AO22X1 U4062 (.IN1(n7013), .IN2(n2780), .IN3(\key_mem[7][30] ), .IN4(n7242), .Q(n4888)
          );
   AO22X1 U4063 (.IN1(n6756), .IN2(n2780), .IN3(\key_mem[8][30] ), .IN4(n6718), .Q(n4889)
          );
   AO22X1 U4064 (.IN1(n7224), .IN2(n2780), .IN3(\key_mem[9][30] ), .IN4(n7214), .Q(n4890)
          );
   AO22X1 U4065 (.IN1(n6803), .IN2(n2780), .IN3(\key_mem[10][30] ), .IN4(n6765), .Q(n4891)
          );
   AO22X1 U4066 (.IN1(n7200), .IN2(n2780), .IN3(\key_mem[11][30] ), .IN4(n7190), .Q(n4892)
          );
   AO22X1 U4067 (.IN1(n6832), .IN2(n2780), .IN3(\key_mem[12][30] ), .IN4(n7184), .Q(n4893)
          );
   AO22X1 U4068 (.IN1(n7179), .IN2(n2780), .IN3(\key_mem[13][30] ), .IN4(n7169), .Q(n4894)
          );
   AO22X1 U4069 (.IN1(n6995), .IN2(n2780), .IN3(\key_mem[14][30] ), .IN4(n7150), .Q(n4895)
          );
   AO221X1 U4070 (.IN1(n7134), .IN2(n2781), .IN3(key[158]), .IN4(n7297), .IN5(n2782), .Q(
          n2780));
   AO222X1 U4071 (.IN1(n7110), .IN2(n2783), .IN3(key[30]), .IN4(n7079), .IN5(n7046), .IN6(
          n2784), .Q(n2782));
   AO22X1 U4072 (.IN1(n7312), .IN2(n2785), .IN3(\key_mem[0][29] ), .IN4(n6930), .Q(n4896)
          );
   AO22X1 U4073 (.IN1(n6927), .IN2(n2785), .IN3(\key_mem[1][29] ), .IN4(n6815), .Q(n4897)
          );
   AO22X1 U4074 (.IN1(n6855), .IN2(n2785), .IN3(\key_mem[2][29] ), .IN4(n6846), .Q(n4898)
          );
   AO22X1 U4075 (.IN1(n6806), .IN2(n2785), .IN3(\key_mem[3][29] ), .IN4(n6863), .Q(n4899)
          );
   AO22X1 U4076 (.IN1(n6921), .IN2(n2785), .IN3(\key_mem[4][29] ), .IN4(n6919), .Q(n4900)
          );
   AO22X1 U4077 (.IN1(n7275), .IN2(n2785), .IN3(\key_mem[5][29] ), .IN4(n7270), .Q(n4901)
          );
   AO22X1 U4078 (.IN1(n7263), .IN2(n2785), .IN3(\key_mem[6][29] ), .IN4(n7253), .Q(n4902)
          );
   AO22X1 U4079 (.IN1(n7014), .IN2(n2785), .IN3(\key_mem[7][29] ), .IN4(n7237), .Q(n4903)
          );
   AO22X1 U4080 (.IN1(n6757), .IN2(n2785), .IN3(\key_mem[8][29] ), .IN4(n6719), .Q(n4904)
          );
   AO22X1 U4081 (.IN1(n7219), .IN2(n2785), .IN3(\key_mem[9][29] ), .IN4(n7214), .Q(n4905)
          );
   AO22X1 U4082 (.IN1(n6804), .IN2(n2785), .IN3(\key_mem[10][29] ), .IN4(n6766), .Q(n4906)
          );
   AO22X1 U4083 (.IN1(n7195), .IN2(n2785), .IN3(\key_mem[11][29] ), .IN4(n7190), .Q(n4907)
          );
   AO22X1 U4084 (.IN1(n6827), .IN2(n2785), .IN3(\key_mem[12][29] ), .IN4(n6985), .Q(n4908)
          );
   AO22X1 U4085 (.IN1(n7174), .IN2(n2785), .IN3(\key_mem[13][29] ), .IN4(n7169), .Q(n4909)
          );
   AO22X1 U4086 (.IN1(n6996), .IN2(n2785), .IN3(\key_mem[14][29] ), .IN4(n7151), .Q(n4910)
          );
   AO221X1 U4087 (.IN1(n7134), .IN2(n2786), .IN3(key[157]), .IN4(n7298), .IN5(n2787), .Q(
          n2785));
   AO222X1 U4088 (.IN1(n7110), .IN2(n2788), .IN3(key[29]), .IN4(n7079), .IN5(n7046), .IN6(
          n2789), .Q(n2787));
   AO22X1 U4089 (.IN1(n2276), .IN2(n2790), .IN3(\key_mem[0][28] ), .IN4(n6930), .Q(n4911)
          );
   AO22X1 U4090 (.IN1(n6809), .IN2(n2790), .IN3(\key_mem[1][28] ), .IN4(n6821), .Q(n4912)
          );
   AO22X1 U4091 (.IN1(n6855), .IN2(n2790), .IN3(\key_mem[2][28] ), .IN4(n6851), .Q(n4913)
          );
   AO22X1 U4092 (.IN1(n6875), .IN2(n2790), .IN3(\key_mem[3][28] ), .IN4(n6865), .Q(n4914)
          );
   AO22X1 U4093 (.IN1(n6888), .IN2(n2790), .IN3(\key_mem[4][28] ), .IN4(n6925), .Q(n4915)
          );
   AO22X1 U4094 (.IN1(n7274), .IN2(n2790), .IN3(\key_mem[5][28] ), .IN4(n7282), .Q(n4916)
          );
   AO22X1 U4095 (.IN1(n6969), .IN2(n2790), .IN3(\key_mem[6][28] ), .IN4(n7258), .Q(n4917)
          );
   AO22X1 U4096 (.IN1(n7013), .IN2(n2790), .IN3(\key_mem[7][28] ), .IN4(n7236), .Q(n4918)
          );
   AO22X1 U4097 (.IN1(n6758), .IN2(n2790), .IN3(\key_mem[8][28] ), .IN4(n6720), .Q(n4919)
          );
   AO22X1 U4098 (.IN1(n7218), .IN2(n2790), .IN3(\key_mem[9][28] ), .IN4(n7226), .Q(n4920)
          );
   AO22X1 U4099 (.IN1(n6805), .IN2(n2790), .IN3(\key_mem[10][28] ), .IN4(n6767), .Q(n4921)
          );
   AO22X1 U4100 (.IN1(n7194), .IN2(n2790), .IN3(\key_mem[11][28] ), .IN4(n7202), .Q(n4922)
          );
   AO22X1 U4101 (.IN1(n6837), .IN2(n2790), .IN3(\key_mem[12][28] ), .IN4(n6830), .Q(n4923)
          );
   AO22X1 U4102 (.IN1(n7173), .IN2(n2790), .IN3(\key_mem[13][28] ), .IN4(n7181), .Q(n4924)
          );
   AO22X1 U4103 (.IN1(n7158), .IN2(n2790), .IN3(\key_mem[14][28] ), .IN4(n7148), .Q(n4925)
          );
   AO221X1 U4104 (.IN1(n7134), .IN2(n2791), .IN3(key[156]), .IN4(n7304), .IN5(n2792), .Q(
          n2790));
   AO222X1 U4105 (.IN1(n7110), .IN2(n2793), .IN3(key[28]), .IN4(n7079), .IN5(n7046), .IN6(
          n2794), .Q(n2792));
   AO22X1 U4106 (.IN1(n7294), .IN2(n2795), .IN3(\key_mem[0][27] ), .IN4(n6930), .Q(n4926)
          );
   AO22X1 U4107 (.IN1(n6812), .IN2(n2795), .IN3(\key_mem[1][27] ), .IN4(n6822), .Q(n4927)
          );
   AO22X1 U4108 (.IN1(n6853), .IN2(n2795), .IN3(\key_mem[2][27] ), .IN4(n6844), .Q(n4928)
          );
   AO22X1 U4109 (.IN1(n6870), .IN2(n2795), .IN3(\key_mem[3][27] ), .IN4(n6865), .Q(n4929)
          );
   AO22X1 U4110 (.IN1(n7287), .IN2(n2795), .IN3(\key_mem[4][27] ), .IN4(n6890), .Q(n4930)
          );
   AO22X1 U4111 (.IN1(n6974), .IN2(n2795), .IN3(\key_mem[5][27] ), .IN4(n7273), .Q(n4931)
          );
   AO22X1 U4112 (.IN1(n7016), .IN2(n2795), .IN3(\key_mem[6][27] ), .IN4(n2283), .Q(n4932)
          );
   AO22X1 U4113 (.IN1(n7013), .IN2(n2795), .IN3(\key_mem[7][27] ), .IN4(n2284), .Q(n4933)
          );
   AO22X1 U4114 (.IN1(n6750), .IN2(n2795), .IN3(\key_mem[8][27] ), .IN4(n6725), .Q(n4934)
          );
   AO22X1 U4115 (.IN1(n6976), .IN2(n2795), .IN3(\key_mem[9][27] ), .IN4(n7217), .Q(n4935)
          );
   AO22X1 U4116 (.IN1(n6797), .IN2(n2795), .IN3(\key_mem[10][27] ), .IN4(n6772), .Q(n4936)
          );
   AO22X1 U4117 (.IN1(n6978), .IN2(n2795), .IN3(\key_mem[11][27] ), .IN4(n7193), .Q(n4937)
          );
   AO22X1 U4118 (.IN1(n7183), .IN2(n2795), .IN3(\key_mem[12][27] ), .IN4(n6830), .Q(n4938)
          );
   AO22X1 U4119 (.IN1(n6980), .IN2(n2795), .IN3(\key_mem[13][27] ), .IN4(n7172), .Q(n4939)
          );
   AO22X1 U4120 (.IN1(n7163), .IN2(n2795), .IN3(\key_mem[14][27] ), .IN4(n7149), .Q(n4940)
          );
   AO221X1 U4121 (.IN1(n7134), .IN2(n2796), .IN3(key[155]), .IN4(n7302), .IN5(n2797), .Q(
          n2795));
   AO222X1 U4122 (.IN1(n7110), .IN2(n2798), .IN3(key[27]), .IN4(n7079), .IN5(n7046), .IN6(
          n2799), .Q(n2797));
   AO22X1 U4123 (.IN1(n7293), .IN2(n2800), .IN3(\key_mem[0][26] ), .IN4(n6930), .Q(n4941)
          );
   AO22X1 U4124 (.IN1(n6808), .IN2(n2800), .IN3(\key_mem[1][26] ), .IN4(n6819), .Q(n4942)
          );
   AO22X1 U4125 (.IN1(n6858), .IN2(n2800), .IN3(\key_mem[2][26] ), .IN4(n6851), .Q(n4943)
          );
   AO22X1 U4126 (.IN1(n6870), .IN2(n2800), .IN3(\key_mem[3][26] ), .IN4(n6863), .Q(n4944)
          );
   AO22X1 U4127 (.IN1(n6889), .IN2(n2800), .IN3(\key_mem[4][26] ), .IN4(n7284), .Q(n4945)
          );
   AO22X1 U4128 (.IN1(n7277), .IN2(n2800), .IN3(\key_mem[5][26] ), .IN4(n7272), .Q(n4946)
          );
   AO22X1 U4129 (.IN1(n7017), .IN2(n2800), .IN3(\key_mem[6][26] ), .IN4(n7015), .Q(n4947)
          );
   AO22X1 U4130 (.IN1(n7248), .IN2(n2800), .IN3(\key_mem[7][26] ), .IN4(n7012), .Q(n4948)
          );
   AO22X1 U4131 (.IN1(n6751), .IN2(n2800), .IN3(\key_mem[8][26] ), .IN4(n6721), .Q(n4949)
          );
   AO22X1 U4132 (.IN1(n7221), .IN2(n2800), .IN3(\key_mem[9][26] ), .IN4(n7216), .Q(n4950)
          );
   AO22X1 U4133 (.IN1(n6798), .IN2(n2800), .IN3(\key_mem[10][26] ), .IN4(n6768), .Q(n4951)
          );
   AO22X1 U4134 (.IN1(n7197), .IN2(n2800), .IN3(\key_mem[11][26] ), .IN4(n7192), .Q(n4952)
          );
   AO22X1 U4135 (.IN1(n6827), .IN2(n2800), .IN3(\key_mem[12][26] ), .IN4(n6981), .Q(n4953)
          );
   AO22X1 U4136 (.IN1(n7176), .IN2(n2800), .IN3(\key_mem[13][26] ), .IN4(n7171), .Q(n4954)
          );
   AO22X1 U4137 (.IN1(n7162), .IN2(n2800), .IN3(\key_mem[14][26] ), .IN4(n7156), .Q(n4955)
          );
   AO221X1 U4138 (.IN1(n7134), .IN2(n2801), .IN3(key[154]), .IN4(n7303), .IN5(n2802), .Q(
          n2800));
   AO222X1 U4139 (.IN1(n7110), .IN2(n2803), .IN3(key[26]), .IN4(n7079), .IN5(n7046), .IN6(
          n2804), .Q(n2802));
   AO22X1 U4140 (.IN1(n7292), .IN2(n2805), .IN3(\key_mem[0][25] ), .IN4(n6930), .Q(n4956)
          );
   AO22X1 U4141 (.IN1(n6812), .IN2(n2805), .IN3(\key_mem[1][25] ), .IN4(n6820), .Q(n4957)
          );
   AO22X1 U4142 (.IN1(n6857), .IN2(n2805), .IN3(\key_mem[2][25] ), .IN4(n6842), .Q(n4958)
          );
   AO22X1 U4143 (.IN1(n6869), .IN2(n2805), .IN3(\key_mem[3][25] ), .IN4(n6862), .Q(n4959)
          );
   AO22X1 U4144 (.IN1(n6990), .IN2(n2805), .IN3(\key_mem[4][25] ), .IN4(n7289), .Q(n4960)
          );
   AO22X1 U4145 (.IN1(n7279), .IN2(n2805), .IN3(\key_mem[5][25] ), .IN4(n2282), .Q(n4961)
          );
   AO22X1 U4146 (.IN1(n7266), .IN2(n2805), .IN3(\key_mem[6][25] ), .IN4(n7257), .Q(n4962)
          );
   AO22X1 U4147 (.IN1(n7014), .IN2(n2805), .IN3(\key_mem[7][25] ), .IN4(n7243), .Q(n4963)
          );
   AO22X1 U4148 (.IN1(n6752), .IN2(n2805), .IN3(\key_mem[8][25] ), .IN4(n6722), .Q(n4964)
          );
   AO22X1 U4149 (.IN1(n7223), .IN2(n2805), .IN3(\key_mem[9][25] ), .IN4(n2286), .Q(n4965)
          );
   AO22X1 U4150 (.IN1(n6799), .IN2(n2805), .IN3(\key_mem[10][25] ), .IN4(n6769), .Q(n4966)
          );
   AO22X1 U4151 (.IN1(n7199), .IN2(n2805), .IN3(\key_mem[11][25] ), .IN4(n2288), .Q(n4967)
          );
   AO22X1 U4152 (.IN1(n6826), .IN2(n2805), .IN3(\key_mem[12][25] ), .IN4(n6839), .Q(n4968)
          );
   AO22X1 U4153 (.IN1(n7178), .IN2(n2805), .IN3(\key_mem[13][25] ), .IN4(n2290), .Q(n4969)
          );
   AO22X1 U4154 (.IN1(n7161), .IN2(n2805), .IN3(\key_mem[14][25] ), .IN4(n7157), .Q(n4970)
          );
   AO221X1 U4155 (.IN1(n7134), .IN2(n2806), .IN3(key[153]), .IN4(n7308), .IN5(n2807), .Q(
          n2805));
   AO222X1 U4156 (.IN1(n7110), .IN2(n2808), .IN3(key[25]), .IN4(n7079), .IN5(n7046), .IN6(
          n2809), .Q(n2807));
   AO22X1 U4157 (.IN1(n7291), .IN2(n2810), .IN3(\key_mem[0][24] ), .IN4(n6930), .Q(n4971)
          );
   AO22X1 U4158 (.IN1(n6813), .IN2(n2810), .IN3(\key_mem[1][24] ), .IN4(n6825), .Q(n4972)
          );
   AO22X1 U4159 (.IN1(n6854), .IN2(n2810), .IN3(\key_mem[2][24] ), .IN4(n6844), .Q(n4973)
          );
   AO22X1 U4160 (.IN1(n6806), .IN2(n2810), .IN3(\key_mem[3][24] ), .IN4(n6862), .Q(n4974)
          );
   AO22X1 U4161 (.IN1(n6889), .IN2(n2810), .IN3(\key_mem[4][24] ), .IN4(n6919), .Q(n4975)
          );
   AO22X1 U4162 (.IN1(n7019), .IN2(n2810), .IN3(\key_mem[5][24] ), .IN4(n7018), .Q(n4976)
          );
   AO22X1 U4163 (.IN1(n7263), .IN2(n2810), .IN3(\key_mem[6][24] ), .IN4(n7015), .Q(n4977)
          );
   AO22X1 U4164 (.IN1(n7244), .IN2(n2810), .IN3(\key_mem[7][24] ), .IN4(n7235), .Q(n4978)
          );
   AO22X1 U4165 (.IN1(n6750), .IN2(n2810), .IN3(\key_mem[8][24] ), .IN4(n6717), .Q(n4979)
          );
   AO22X1 U4166 (.IN1(n7008), .IN2(n2810), .IN3(\key_mem[9][24] ), .IN4(n7007), .Q(n4980)
          );
   AO22X1 U4167 (.IN1(n6797), .IN2(n2810), .IN3(\key_mem[10][24] ), .IN4(n6764), .Q(n4981)
          );
   AO22X1 U4168 (.IN1(n7003), .IN2(n2810), .IN3(\key_mem[11][24] ), .IN4(n7002), .Q(n4982)
          );
   AO22X1 U4169 (.IN1(n6835), .IN2(n2810), .IN3(\key_mem[12][24] ), .IN4(n6828), .Q(n4983)
          );
   AO22X1 U4170 (.IN1(n6998), .IN2(n2810), .IN3(\key_mem[13][24] ), .IN4(n6997), .Q(n4984)
          );
   AO22X1 U4171 (.IN1(n6995), .IN2(n2810), .IN3(\key_mem[14][24] ), .IN4(n7154), .Q(n4985)
          );
   AO221X1 U4172 (.IN1(n7134), .IN2(n2811), .IN3(key[152]), .IN4(n7295), .IN5(n2812), .Q(
          n2810));
   AO222X1 U4173 (.IN1(n7110), .IN2(n2813), .IN3(key[24]), .IN4(n7079), .IN5(n7046), .IN6(
          n2814), .Q(n2812));
   AO22X1 U4174 (.IN1(n7290), .IN2(n2815), .IN3(\key_mem[0][23] ), .IN4(n6929), .Q(n4986)
          );
   AO22X1 U4175 (.IN1(n6926), .IN2(n2815), .IN3(\key_mem[1][23] ), .IN4(n6822), .Q(n4987)
          );
   AO22X1 U4176 (.IN1(n6855), .IN2(n2815), .IN3(\key_mem[2][23] ), .IN4(n6843), .Q(n4988)
          );
   AO22X1 U4177 (.IN1(n6871), .IN2(n2815), .IN3(\key_mem[3][23] ), .IN4(n6876), .Q(n4989)
          );
   AO22X1 U4178 (.IN1(n7288), .IN2(n2815), .IN3(\key_mem[4][23] ), .IN4(n6917), .Q(n4990)
          );
   AO22X1 U4179 (.IN1(n6973), .IN2(n2815), .IN3(\key_mem[5][23] ), .IN4(n7018), .Q(n4991)
          );
   AO22X1 U4180 (.IN1(n7016), .IN2(n2815), .IN3(\key_mem[6][23] ), .IN4(n2283), .Q(n4992)
          );
   AO22X1 U4181 (.IN1(n7245), .IN2(n2815), .IN3(\key_mem[7][23] ), .IN4(n7236), .Q(n4993)
          );
   AO22X1 U4182 (.IN1(n6754), .IN2(n2815), .IN3(\key_mem[8][23] ), .IN4(n6746), .Q(n4994)
          );
   AO22X1 U4183 (.IN1(n6975), .IN2(n2815), .IN3(\key_mem[9][23] ), .IN4(n7007), .Q(n4995)
          );
   AO22X1 U4184 (.IN1(n6801), .IN2(n2815), .IN3(\key_mem[10][23] ), .IN4(n6793), .Q(n4996)
          );
   AO22X1 U4185 (.IN1(n6977), .IN2(n2815), .IN3(\key_mem[11][23] ), .IN4(n7002), .Q(n4997)
          );
   AO22X1 U4186 (.IN1(n6835), .IN2(n2815), .IN3(\key_mem[12][23] ), .IN4(n6828), .Q(n4998)
          );
   AO22X1 U4187 (.IN1(n6979), .IN2(n2815), .IN3(\key_mem[13][23] ), .IN4(n6997), .Q(n4999)
          );
   AO22X1 U4188 (.IN1(n6971), .IN2(n2815), .IN3(\key_mem[14][23] ), .IN4(n7155), .Q(n5000)
          );
   AO221X1 U4189 (.IN1(n7134), .IN2(n2816), .IN3(key[151]), .IN4(n7304), .IN5(n2817), .Q(
          n2815));
   AO222X1 U4190 (.IN1(n7110), .IN2(n2818), .IN3(key[23]), .IN4(n7079), .IN5(n7046), .IN6(
          n2819), .Q(n2817));
   AO22X1 U4191 (.IN1(n7299), .IN2(n2820), .IN3(\key_mem[0][22] ), .IN4(n6929), .Q(n5001)
          );
   AO22X1 U4192 (.IN1(n6811), .IN2(n2820), .IN3(\key_mem[1][22] ), .IN4(n6823), .Q(n5002)
          );
   AO22X1 U4193 (.IN1(n6856), .IN2(n2820), .IN3(\key_mem[2][22] ), .IN4(n6844), .Q(n5003)
          );
   AO22X1 U4194 (.IN1(n6806), .IN2(n2820), .IN3(\key_mem[3][22] ), .IN4(n6864), .Q(n5004)
          );
   AO22X1 U4195 (.IN1(n6889), .IN2(n2820), .IN3(\key_mem[4][22] ), .IN4(n6918), .Q(n5005)
          );
   AO22X1 U4196 (.IN1(n7019), .IN2(n2820), .IN3(\key_mem[5][22] ), .IN4(n7273), .Q(n5006)
          );
   AO22X1 U4197 (.IN1(n7017), .IN2(n2820), .IN3(\key_mem[6][22] ), .IN4(n7255), .Q(n5007)
          );
   AO22X1 U4198 (.IN1(n7246), .IN2(n2820), .IN3(\key_mem[7][22] ), .IN4(n7237), .Q(n5008)
          );
   AO22X1 U4199 (.IN1(n6755), .IN2(n2820), .IN3(\key_mem[8][22] ), .IN4(n6745), .Q(n5009)
          );
   AO22X1 U4200 (.IN1(n7008), .IN2(n2820), .IN3(\key_mem[9][22] ), .IN4(n7217), .Q(n5010)
          );
   AO22X1 U4201 (.IN1(n6802), .IN2(n2820), .IN3(\key_mem[10][22] ), .IN4(n6792), .Q(n5011)
          );
   AO22X1 U4202 (.IN1(n7003), .IN2(n2820), .IN3(\key_mem[11][22] ), .IN4(n7193), .Q(n5012)
          );
   AO22X1 U4203 (.IN1(n6829), .IN2(n2820), .IN3(\key_mem[12][22] ), .IN4(n6836), .Q(n5013)
          );
   AO22X1 U4204 (.IN1(n6998), .IN2(n2820), .IN3(\key_mem[13][22] ), .IN4(n7172), .Q(n5014)
          );
   AO22X1 U4205 (.IN1(n7162), .IN2(n2820), .IN3(\key_mem[14][22] ), .IN4(n7165), .Q(n5015)
          );
   AO221X1 U4206 (.IN1(n7134), .IN2(n2821), .IN3(key[150]), .IN4(n7308), .IN5(n2822), .Q(
          n2820));
   AO222X1 U4207 (.IN1(n7110), .IN2(n2823), .IN3(key[22]), .IN4(n7079), .IN5(n7046), .IN6(
          n2824), .Q(n2822));
   AO22X1 U4208 (.IN1(n7298), .IN2(n2825), .IN3(\key_mem[0][21] ), .IN4(n6929), .Q(n5016)
          );
   AO22X1 U4209 (.IN1(n6810), .IN2(n2825), .IN3(\key_mem[1][21] ), .IN4(n6824), .Q(n5017)
          );
   AO22X1 U4210 (.IN1(n6856), .IN2(n2825), .IN3(\key_mem[2][21] ), .IN4(n6851), .Q(n5018)
          );
   AO22X1 U4211 (.IN1(n6870), .IN2(n2825), .IN3(\key_mem[3][21] ), .IN4(n6864), .Q(n5019)
          );
   AO22X1 U4212 (.IN1(n7022), .IN2(n2825), .IN3(\key_mem[4][21] ), .IN4(n6915), .Q(n5020)
          );
   AO22X1 U4213 (.IN1(n7278), .IN2(n2825), .IN3(\key_mem[5][21] ), .IN4(n2282), .Q(n5021)
          );
   AO22X1 U4214 (.IN1(n6970), .IN2(n2825), .IN3(\key_mem[6][21] ), .IN4(n7258), .Q(n5022)
          );
   AO22X1 U4215 (.IN1(n7247), .IN2(n2825), .IN3(\key_mem[7][21] ), .IN4(n7243), .Q(n5023)
          );
   AO22X1 U4216 (.IN1(n6756), .IN2(n2825), .IN3(\key_mem[8][21] ), .IN4(n6743), .Q(n5024)
          );
   AO22X1 U4217 (.IN1(n7222), .IN2(n2825), .IN3(\key_mem[9][21] ), .IN4(n2286), .Q(n5025)
          );
   AO22X1 U4218 (.IN1(n6803), .IN2(n2825), .IN3(\key_mem[10][21] ), .IN4(n6790), .Q(n5026)
          );
   AO22X1 U4219 (.IN1(n7198), .IN2(n2825), .IN3(\key_mem[11][21] ), .IN4(n2288), .Q(n5027)
          );
   AO22X1 U4220 (.IN1(n7183), .IN2(n2825), .IN3(\key_mem[12][21] ), .IN4(n6982), .Q(n5028)
          );
   AO22X1 U4221 (.IN1(n7177), .IN2(n2825), .IN3(\key_mem[13][21] ), .IN4(n2290), .Q(n5029)
          );
   AO22X1 U4222 (.IN1(n6995), .IN2(n2825), .IN3(\key_mem[14][21] ), .IN4(n7148), .Q(n5030)
          );
   AO221X1 U4223 (.IN1(n7134), .IN2(n2826), .IN3(key[149]), .IN4(n7306), .IN5(n2827), .Q(
          n2825));
   AO222X1 U4224 (.IN1(n7110), .IN2(n2828), .IN3(key[21]), .IN4(n7079), .IN5(n7046), .IN6(
          n2829), .Q(n2827));
   AO22X1 U4225 (.IN1(n7306), .IN2(n2830), .IN3(\key_mem[0][20] ), .IN4(n6929), .Q(n5031)
          );
   AO22X1 U4226 (.IN1(n6810), .IN2(n2830), .IN3(\key_mem[1][20] ), .IN4(n6825), .Q(n5032)
          );
   AO22X1 U4227 (.IN1(n6856), .IN2(n2830), .IN3(\key_mem[2][20] ), .IN4(n6847), .Q(n5033)
          );
   AO22X1 U4228 (.IN1(n6869), .IN2(n2830), .IN3(\key_mem[3][20] ), .IN4(n6863), .Q(n5034)
          );
   AO22X1 U4229 (.IN1(n6888), .IN2(n2830), .IN3(\key_mem[4][20] ), .IN4(n7285), .Q(n5035)
          );
   AO22X1 U4230 (.IN1(n7275), .IN2(n2830), .IN3(\key_mem[5][20] ), .IN4(n7269), .Q(n5036)
          );
   AO22X1 U4231 (.IN1(n6970), .IN2(n2830), .IN3(\key_mem[6][20] ), .IN4(n7252), .Q(n5037)
          );
   AO22X1 U4232 (.IN1(n7248), .IN2(n2830), .IN3(\key_mem[7][20] ), .IN4(n7239), .Q(n5038)
          );
   AO22X1 U4233 (.IN1(n6755), .IN2(n2830), .IN3(\key_mem[8][20] ), .IN4(n6742), .Q(n5039)
          );
   AO22X1 U4234 (.IN1(n7219), .IN2(n2830), .IN3(\key_mem[9][20] ), .IN4(n7214), .Q(n5040)
          );
   AO22X1 U4235 (.IN1(n6802), .IN2(n2830), .IN3(\key_mem[10][20] ), .IN4(n6789), .Q(n5041)
          );
   AO22X1 U4236 (.IN1(n7195), .IN2(n2830), .IN3(\key_mem[11][20] ), .IN4(n7190), .Q(n5042)
          );
   AO22X1 U4237 (.IN1(n7001), .IN2(n2830), .IN3(\key_mem[12][20] ), .IN4(n6838), .Q(n5043)
          );
   AO22X1 U4238 (.IN1(n7174), .IN2(n2830), .IN3(\key_mem[13][20] ), .IN4(n7169), .Q(n5044)
          );
   AO22X1 U4239 (.IN1(n6996), .IN2(n2830), .IN3(\key_mem[14][20] ), .IN4(n7154), .Q(n5045)
          );
   AO221X1 U4240 (.IN1(n7134), .IN2(n2831), .IN3(key[148]), .IN4(n7300), .IN5(n2832), .Q(
          n2830));
   AO222X1 U4241 (.IN1(n7110), .IN2(n2833), .IN3(key[20]), .IN4(n7079), .IN5(n7046), .IN6(
          n2834), .Q(n2832));
   AO22X1 U4242 (.IN1(n7303), .IN2(n2835), .IN3(\key_mem[0][19] ), .IN4(n6929), .Q(n5046)
          );
   AO22X1 U4243 (.IN1(n6808), .IN2(n2835), .IN3(\key_mem[1][19] ), .IN4(n6814), .Q(n5047)
          );
   AO22X1 U4244 (.IN1(n6854), .IN2(n2835), .IN3(\key_mem[2][19] ), .IN4(n6848), .Q(n5048)
          );
   AO22X1 U4245 (.IN1(n6873), .IN2(n2835), .IN3(\key_mem[3][19] ), .IN4(n6877), .Q(n5049)
          );
   AO22X1 U4246 (.IN1(n7287), .IN2(n2835), .IN3(\key_mem[4][19] ), .IN4(n6923), .Q(n5050)
          );
   AO22X1 U4247 (.IN1(n7275), .IN2(n2835), .IN3(\key_mem[5][19] ), .IN4(n7273), .Q(n5051)
          );
   AO22X1 U4248 (.IN1(n6970), .IN2(n2835), .IN3(\key_mem[6][19] ), .IN4(n2283), .Q(n5052)
          );
   AO22X1 U4249 (.IN1(n7014), .IN2(n2835), .IN3(\key_mem[7][19] ), .IN4(n7237), .Q(n5053)
          );
   AO22X1 U4250 (.IN1(n6756), .IN2(n2835), .IN3(\key_mem[8][19] ), .IN4(n6716), .Q(n5054)
          );
   AO22X1 U4251 (.IN1(n7219), .IN2(n2835), .IN3(\key_mem[9][19] ), .IN4(n7211), .Q(n5055)
          );
   AO22X1 U4252 (.IN1(n6803), .IN2(n2835), .IN3(\key_mem[10][19] ), .IN4(n6763), .Q(n5056)
          );
   AO22X1 U4253 (.IN1(n7195), .IN2(n2835), .IN3(\key_mem[11][19] ), .IN4(n7187), .Q(n5057)
          );
   AO22X1 U4254 (.IN1(n6831), .IN2(n2835), .IN3(\key_mem[12][19] ), .IN4(n6985), .Q(n5058)
          );
   AO22X1 U4255 (.IN1(n7174), .IN2(n2835), .IN3(\key_mem[13][19] ), .IN4(n7166), .Q(n5059)
          );
   AO22X1 U4256 (.IN1(n7159), .IN2(n2835), .IN3(\key_mem[14][19] ), .IN4(n7149), .Q(n5060)
          );
   AO221X1 U4257 (.IN1(n7135), .IN2(n2836), .IN3(key[147]), .IN4(n7298), .IN5(n2837), .Q(
          n2835));
   AO222X1 U4258 (.IN1(n7110), .IN2(n2838), .IN3(key[19]), .IN4(n7080), .IN5(n7047), .IN6(
          n2839), .Q(n2837));
   AO22X1 U4259 (.IN1(n2276), .IN2(n2840), .IN3(\key_mem[0][18] ), .IN4(n6929), .Q(n5061)
          );
   AO22X1 U4260 (.IN1(n6812), .IN2(n2840), .IN3(\key_mem[1][18] ), .IN4(n6825), .Q(n5062)
          );
   AO22X1 U4261 (.IN1(n6855), .IN2(n2840), .IN3(\key_mem[2][18] ), .IN4(n6850), .Q(n5063)
          );
   AO22X1 U4262 (.IN1(n6869), .IN2(n2840), .IN3(\key_mem[3][18] ), .IN4(n6862), .Q(n5064)
          );
   AO22X1 U4263 (.IN1(n6920), .IN2(n2840), .IN3(\key_mem[4][18] ), .IN4(n7284), .Q(n5065)
          );
   AO22X1 U4264 (.IN1(n7274), .IN2(n2840), .IN3(\key_mem[5][18] ), .IN4(n7267), .Q(n5066)
          );
   AO22X1 U4265 (.IN1(n7262), .IN2(n2840), .IN3(\key_mem[6][18] ), .IN4(n7251), .Q(n5067)
          );
   AO22X1 U4266 (.IN1(n7014), .IN2(n2840), .IN3(\key_mem[7][18] ), .IN4(n7240), .Q(n5068)
          );
   AO22X1 U4267 (.IN1(n6758), .IN2(n2840), .IN3(\key_mem[8][18] ), .IN4(n6715), .Q(n5069)
          );
   AO22X1 U4268 (.IN1(n7218), .IN2(n2840), .IN3(\key_mem[9][18] ), .IN4(n7211), .Q(n5070)
          );
   AO22X1 U4269 (.IN1(n6805), .IN2(n2840), .IN3(\key_mem[10][18] ), .IN4(n6762), .Q(n5071)
          );
   AO22X1 U4270 (.IN1(n7194), .IN2(n2840), .IN3(\key_mem[11][18] ), .IN4(n7187), .Q(n5072)
          );
   AO22X1 U4271 (.IN1(n6837), .IN2(n2840), .IN3(\key_mem[12][18] ), .IN4(n6834), .Q(n5073)
          );
   AO22X1 U4272 (.IN1(n7173), .IN2(n2840), .IN3(\key_mem[13][18] ), .IN4(n7166), .Q(n5074)
          );
   AO22X1 U4273 (.IN1(n7158), .IN2(n2840), .IN3(\key_mem[14][18] ), .IN4(n7156), .Q(n5075)
          );
   AO222X1 U4275 (.IN1(n7110), .IN2(n2843), .IN3(key[18]), .IN4(n7080), .IN5(n7047), .IN6(
          n2844), .Q(n2842));
   AO22X1 U4276 (.IN1(n7292), .IN2(n2845), .IN3(\key_mem[0][17] ), .IN4(n6929), .Q(n5076)
          );
   AO22X1 U4277 (.IN1(n6927), .IN2(n2845), .IN3(\key_mem[1][17] ), .IN4(n6814), .Q(n5077)
          );
   AO22X1 U4278 (.IN1(n6856), .IN2(n2845), .IN3(\key_mem[2][17] ), .IN4(n6844), .Q(n5078)
          );
   AO22X1 U4279 (.IN1(n6989), .IN2(n2845), .IN3(\key_mem[3][17] ), .IN4(n6867), .Q(n5079)
          );
   AO22X1 U4280 (.IN1(n7288), .IN2(n2845), .IN3(\key_mem[4][17] ), .IN4(n7289), .Q(n5080)
          );
   AO22X1 U4281 (.IN1(n7276), .IN2(n2845), .IN3(\key_mem[5][17] ), .IN4(n7271), .Q(n5081)
          );
   AO22X1 U4282 (.IN1(n7264), .IN2(n2845), .IN3(\key_mem[6][17] ), .IN4(n7259), .Q(n5082)
          );
   AO22X1 U4283 (.IN1(n7250), .IN2(n2845), .IN3(\key_mem[7][17] ), .IN4(n7238), .Q(n5083)
          );
   AO22X1 U4284 (.IN1(n6751), .IN2(n2845), .IN3(\key_mem[8][17] ), .IN4(n6719), .Q(n5084)
          );
   AO22X1 U4285 (.IN1(n7220), .IN2(n2845), .IN3(\key_mem[9][17] ), .IN4(n7214), .Q(n5085)
          );
   AO22X1 U4286 (.IN1(n6798), .IN2(n2845), .IN3(\key_mem[10][17] ), .IN4(n6766), .Q(n5086)
          );
   AO22X1 U4287 (.IN1(n7196), .IN2(n2845), .IN3(\key_mem[11][17] ), .IN4(n7190), .Q(n5087)
          );
   AO22X1 U4288 (.IN1(n6987), .IN2(n2845), .IN3(\key_mem[12][17] ), .IN4(n6984), .Q(n5088)
          );
   AO22X1 U4289 (.IN1(n7175), .IN2(n2845), .IN3(\key_mem[13][17] ), .IN4(n7169), .Q(n5089)
          );
   AO22X1 U4290 (.IN1(n7162), .IN2(n2845), .IN3(\key_mem[14][17] ), .IN4(n7157), .Q(n5090)
          );
   AO221X1 U4291 (.IN1(n7135), .IN2(n2846), .IN3(key[145]), .IN4(n7307), .IN5(n2847), .Q(
          n2845));
   AO222X1 U4292 (.IN1(n7109), .IN2(n2848), .IN3(key[17]), .IN4(n7080), .IN5(n7047), .IN6(
          n2849), .Q(n2847));
   AO22X1 U4293 (.IN1(n7291), .IN2(n2850), .IN3(\key_mem[0][16] ), .IN4(n6929), .Q(n5091)
          );
   AO22X1 U4294 (.IN1(n6811), .IN2(n2850), .IN3(\key_mem[1][16] ), .IN4(n6815), .Q(n5092)
          );
   AO22X1 U4295 (.IN1(n6988), .IN2(n2850), .IN3(\key_mem[2][16] ), .IN4(n6848), .Q(n5093)
          );
   AO22X1 U4296 (.IN1(n6989), .IN2(n2850), .IN3(\key_mem[3][16] ), .IN4(n6860), .Q(n5094)
          );
   AO22X1 U4297 (.IN1(n6886), .IN2(n2850), .IN3(\key_mem[4][16] ), .IN4(n7021), .Q(n5095)
          );
   AO22X1 U4298 (.IN1(n7277), .IN2(n2850), .IN3(\key_mem[5][16] ), .IN4(n2282), .Q(n5096)
          );
   AO22X1 U4299 (.IN1(n7263), .IN2(n2850), .IN3(\key_mem[6][16] ), .IN4(n7258), .Q(n5097)
          );
   AO22X1 U4300 (.IN1(n7244), .IN2(n2850), .IN3(\key_mem[7][16] ), .IN4(n7239), .Q(n5098)
          );
   AO22X1 U4301 (.IN1(n6748), .IN2(n2850), .IN3(\key_mem[8][16] ), .IN4(n6714), .Q(n5099)
          );
   AO22X1 U4302 (.IN1(n7221), .IN2(n2850), .IN3(\key_mem[9][16] ), .IN4(n2286), .Q(n5100)
          );
   AO22X1 U4303 (.IN1(n6795), .IN2(n2850), .IN3(\key_mem[10][16] ), .IN4(n6761), .Q(n5101)
          );
   AO22X1 U4304 (.IN1(n7197), .IN2(n2850), .IN3(\key_mem[11][16] ), .IN4(n2288), .Q(n5102)
          );
   AO22X1 U4305 (.IN1(n6826), .IN2(n2850), .IN3(\key_mem[12][16] ), .IN4(n6830), .Q(n5103)
          );
   AO22X1 U4306 (.IN1(n7176), .IN2(n2850), .IN3(\key_mem[13][16] ), .IN4(n2290), .Q(n5104)
          );
   AO22X1 U4307 (.IN1(n7160), .IN2(n2850), .IN3(\key_mem[14][16] ), .IN4(n7154), .Q(n5105)
          );
   AO221X1 U4308 (.IN1(n7135), .IN2(n2851), .IN3(key[144]), .IN4(n7305), .IN5(n2852), .Q(
          n2850));
   AO222X1 U4309 (.IN1(n7109), .IN2(n2853), .IN3(key[16]), .IN4(n7080), .IN5(n7047), .IN6(
          n2854), .Q(n2852));
   AO22X1 U4310 (.IN1(n7290), .IN2(n2855), .IN3(\key_mem[0][15] ), .IN4(n6929), .Q(n5106)
          );
   AO22X1 U4311 (.IN1(n6808), .IN2(n2855), .IN3(\key_mem[1][15] ), .IN4(n6820), .Q(n5107)
          );
   AO22X1 U4312 (.IN1(n6988), .IN2(n2855), .IN3(\key_mem[2][15] ), .IN4(n6843), .Q(n5108)
          );
   AO22X1 U4313 (.IN1(n6873), .IN2(n2855), .IN3(\key_mem[3][15] ), .IN4(n6868), .Q(n5109)
          );
   AO22X1 U4314 (.IN1(n7287), .IN2(n2855), .IN3(\key_mem[4][15] ), .IN4(n6914), .Q(n5110)
          );
   AO22X1 U4315 (.IN1(n6973), .IN2(n2855), .IN3(\key_mem[5][15] ), .IN4(n7271), .Q(n5111)
          );
   AO22X1 U4316 (.IN1(n7262), .IN2(n2855), .IN3(\key_mem[6][15] ), .IN4(n7256), .Q(n5112)
          );
   AO22X1 U4317 (.IN1(n7250), .IN2(n2855), .IN3(\key_mem[7][15] ), .IN4(n7240), .Q(n5113)
          );
   AO22X1 U4318 (.IN1(n6748), .IN2(n2855), .IN3(\key_mem[8][15] ), .IN4(n6714), .Q(n5114)
          );
   AO22X1 U4319 (.IN1(n6975), .IN2(n2855), .IN3(\key_mem[9][15] ), .IN4(n7215), .Q(n5115)
          );
   AO22X1 U4320 (.IN1(n6795), .IN2(n2855), .IN3(\key_mem[10][15] ), .IN4(n6761), .Q(n5116)
          );
   AO22X1 U4321 (.IN1(n6977), .IN2(n2855), .IN3(\key_mem[11][15] ), .IN4(n7191), .Q(n5117)
          );
   AO22X1 U4322 (.IN1(n7001), .IN2(n2855), .IN3(\key_mem[12][15] ), .IN4(n2289), .Q(n5118)
          );
   AO22X1 U4323 (.IN1(n6979), .IN2(n2855), .IN3(\key_mem[13][15] ), .IN4(n7170), .Q(n5119)
          );
   AO22X1 U4324 (.IN1(n6972), .IN2(n2855), .IN3(\key_mem[14][15] ), .IN4(n7155), .Q(n5120)
          );
   AO221X1 U4325 (.IN1(n7135), .IN2(n2856), .IN3(key[143]), .IN4(n7311), .IN5(n2857), .Q(
          n2855));
   AO222X1 U4326 (.IN1(n7109), .IN2(n2858), .IN3(key[15]), .IN4(n7080), .IN5(n7047), .IN6(
          n2859), .Q(n2857));
   AO22X1 U4327 (.IN1(n7299), .IN2(n2860), .IN3(\key_mem[0][14] ), .IN4(n6929), .Q(n5121)
          );
   AO22X1 U4328 (.IN1(n6813), .IN2(n2860), .IN3(\key_mem[1][14] ), .IN4(n6824), .Q(n5122)
          );
   AO22X1 U4329 (.IN1(n6855), .IN2(n2860), .IN3(\key_mem[2][14] ), .IN4(n6846), .Q(n5123)
          );
   AO22X1 U4330 (.IN1(n6989), .IN2(n2860), .IN3(\key_mem[3][14] ), .IN4(n6868), .Q(n5124)
          );
   AO22X1 U4331 (.IN1(n6889), .IN2(n2860), .IN3(\key_mem[4][14] ), .IN4(n6918), .Q(n5125)
          );
   AO22X1 U4332 (.IN1(n6974), .IN2(n2860), .IN3(\key_mem[5][14] ), .IN4(n7272), .Q(n5126)
          );
   AO22X1 U4333 (.IN1(n7261), .IN2(n2860), .IN3(\key_mem[6][14] ), .IN4(n7257), .Q(n5127)
          );
   AO22X1 U4334 (.IN1(n7249), .IN2(n2860), .IN3(\key_mem[7][14] ), .IN4(n7241), .Q(n5128)
          );
   AO22X1 U4335 (.IN1(n6749), .IN2(n2860), .IN3(\key_mem[8][14] ), .IN4(n6719), .Q(n5129)
          );
   AO22X1 U4336 (.IN1(n6976), .IN2(n2860), .IN3(\key_mem[9][14] ), .IN4(n7216), .Q(n5130)
          );
   AO22X1 U4337 (.IN1(n6796), .IN2(n2860), .IN3(\key_mem[10][14] ), .IN4(n6766), .Q(n5131)
          );
   AO22X1 U4338 (.IN1(n6978), .IN2(n2860), .IN3(\key_mem[11][14] ), .IN4(n7192), .Q(n5132)
          );
   AO22X1 U4339 (.IN1(n6829), .IN2(n2860), .IN3(\key_mem[12][14] ), .IN4(n6836), .Q(n5133)
          );
   AO22X1 U4340 (.IN1(n6980), .IN2(n2860), .IN3(\key_mem[13][14] ), .IN4(n7171), .Q(n5134)
          );
   AO22X1 U4341 (.IN1(n7164), .IN2(n2860), .IN3(\key_mem[14][14] ), .IN4(n7147), .Q(n5135)
          );
   AO221X1 U4342 (.IN1(n7135), .IN2(n2861), .IN3(key[142]), .IN4(n7302), .IN5(n2862), .Q(
          n2860));
   AO222X1 U4343 (.IN1(n7109), .IN2(n2863), .IN3(key[14]), .IN4(n7080), .IN5(n7047), .IN6(
          n2864), .Q(n2862));
   AO22X1 U4344 (.IN1(n7298), .IN2(n2865), .IN3(\key_mem[0][13] ), .IN4(n6929), .Q(n5136)
          );
   AO22X1 U4345 (.IN1(n6810), .IN2(n2865), .IN3(\key_mem[1][13] ), .IN4(n6820), .Q(n5137)
          );
   AO22X1 U4346 (.IN1(n6852), .IN2(n2865), .IN3(\key_mem[2][13] ), .IN4(n6843), .Q(n5138)
          );
   AO22X1 U4347 (.IN1(n6872), .IN2(n2865), .IN3(\key_mem[3][13] ), .IN4(n6866), .Q(n5139)
          );
   AO22X1 U4348 (.IN1(n6922), .IN2(n2865), .IN3(\key_mem[4][13] ), .IN4(n7284), .Q(n5140)
          );
   AO22X1 U4349 (.IN1(n6973), .IN2(n2865), .IN3(\key_mem[5][13] ), .IN4(n7282), .Q(n5141)
          );
   AO22X1 U4350 (.IN1(n7262), .IN2(n2865), .IN3(\key_mem[6][13] ), .IN4(n7254), .Q(n5142)
          );
   AO22X1 U4351 (.IN1(n7013), .IN2(n2865), .IN3(\key_mem[7][13] ), .IN4(n7242), .Q(n5143)
          );
   AO22X1 U4352 (.IN1(n6756), .IN2(n2865), .IN3(\key_mem[8][13] ), .IN4(n6717), .Q(n5144)
          );
   AO22X1 U4353 (.IN1(n6975), .IN2(n2865), .IN3(\key_mem[9][13] ), .IN4(n7226), .Q(n5145)
          );
   AO22X1 U4354 (.IN1(n6803), .IN2(n2865), .IN3(\key_mem[10][13] ), .IN4(n6764), .Q(n5146)
          );
   AO22X1 U4355 (.IN1(n6977), .IN2(n2865), .IN3(\key_mem[11][13] ), .IN4(n7202), .Q(n5147)
          );
   AO22X1 U4356 (.IN1(n6840), .IN2(n2865), .IN3(\key_mem[12][13] ), .IN4(n6834), .Q(n5148)
          );
   AO22X1 U4357 (.IN1(n6979), .IN2(n2865), .IN3(\key_mem[13][13] ), .IN4(n7181), .Q(n5149)
          );
   AO22X1 U4358 (.IN1(n7163), .IN2(n2865), .IN3(\key_mem[14][13] ), .IN4(n7165), .Q(n5150)
          );
   AO222X1 U4360 (.IN1(n7109), .IN2(n2868), .IN3(key[13]), .IN4(n7080), .IN5(n7047), .IN6(
          n2869), .Q(n2867));
   AO22X1 U4361 (.IN1(n7297), .IN2(n2870), .IN3(\key_mem[0][12] ), .IN4(n6929), .Q(n5151)
          );
   AO22X1 U4362 (.IN1(n6812), .IN2(n2870), .IN3(\key_mem[1][12] ), .IN4(n6822), .Q(n5152)
          );
   AO22X1 U4363 (.IN1(n6988), .IN2(n2870), .IN3(\key_mem[2][12] ), .IN4(n6850), .Q(n5153)
          );
   AO22X1 U4364 (.IN1(n6871), .IN2(n2870), .IN3(\key_mem[3][12] ), .IN4(n6877), .Q(n5154)
          );
   AO22X1 U4365 (.IN1(n6920), .IN2(n2870), .IN3(\key_mem[4][12] ), .IN4(n6923), .Q(n5155)
          );
   AO22X1 U4366 (.IN1(n7020), .IN2(n2870), .IN3(\key_mem[5][12] ), .IN4(n7267), .Q(n5156)
          );
   AO22X1 U4367 (.IN1(n7266), .IN2(n2870), .IN3(\key_mem[6][12] ), .IN4(n7255), .Q(n5157)
          );
   AO22X1 U4368 (.IN1(n7014), .IN2(n2870), .IN3(\key_mem[7][12] ), .IN4(n7241), .Q(n5158)
          );
   AO22X1 U4369 (.IN1(n6749), .IN2(n2870), .IN3(\key_mem[8][12] ), .IN4(n7228), .Q(n5159)
          );
   AO22X1 U4370 (.IN1(n7009), .IN2(n2870), .IN3(\key_mem[9][12] ), .IN4(n7211), .Q(n5160)
          );
   AO22X1 U4371 (.IN1(n6796), .IN2(n2870), .IN3(\key_mem[10][12] ), .IN4(n7204), .Q(n5161)
          );
   AO22X1 U4372 (.IN1(n7004), .IN2(n2870), .IN3(\key_mem[11][12] ), .IN4(n7187), .Q(n5162)
          );
   AO22X1 U4373 (.IN1(n7001), .IN2(n2870), .IN3(\key_mem[12][12] ), .IN4(n6836), .Q(n5163)
          );
   AO22X1 U4374 (.IN1(n6999), .IN2(n2870), .IN3(\key_mem[13][12] ), .IN4(n7166), .Q(n5164)
          );
   AO22X1 U4375 (.IN1(n6996), .IN2(n2870), .IN3(\key_mem[14][12] ), .IN4(n7147), .Q(n5165)
          );
   AO221X1 U4376 (.IN1(n7135), .IN2(n2871), .IN3(key[140]), .IN4(n7293), .IN5(n2872), .Q(
          n2870));
   AO222X1 U4377 (.IN1(n7109), .IN2(n2873), .IN3(key[12]), .IN4(n7080), .IN5(n7047), .IN6(
          n2874), .Q(n2872));
   AO22X1 U4378 (.IN1(n7296), .IN2(n2875), .IN3(\key_mem[0][11] ), .IN4(n6928), .Q(n5166)
          );
   AO22X1 U4379 (.IN1(n6810), .IN2(n2875), .IN3(\key_mem[1][11] ), .IN4(n6823), .Q(n5167)
          );
   AO22X1 U4380 (.IN1(n6852), .IN2(n2875), .IN3(\key_mem[2][11] ), .IN4(n6846), .Q(n5168)
          );
   AO22X1 U4381 (.IN1(n6806), .IN2(n2875), .IN3(\key_mem[3][11] ), .IN4(n6864), .Q(n5169)
          );
   AO22X1 U4382 (.IN1(n7022), .IN2(n2875), .IN3(\key_mem[4][11] ), .IN4(n6890), .Q(n5170)
          );
   AO22X1 U4383 (.IN1(n7283), .IN2(n2875), .IN3(\key_mem[5][11] ), .IN4(n7271), .Q(n5171)
          );
   AO22X1 U4384 (.IN1(n7264), .IN2(n2875), .IN3(\key_mem[6][11] ), .IN4(n7254), .Q(n5172)
          );
   AO22X1 U4385 (.IN1(n7244), .IN2(n2875), .IN3(\key_mem[7][11] ), .IN4(n7240), .Q(n5173)
          );
   AO22X1 U4386 (.IN1(n6748), .IN2(n2875), .IN3(\key_mem[8][11] ), .IN4(n6734), .Q(n5174)
          );
   AO22X1 U4387 (.IN1(n7227), .IN2(n2875), .IN3(\key_mem[9][11] ), .IN4(n7215), .Q(n5175)
          );
   AO22X1 U4388 (.IN1(n6795), .IN2(n2875), .IN3(\key_mem[10][11] ), .IN4(n6781), .Q(n5176)
          );
   AO22X1 U4389 (.IN1(n7203), .IN2(n2875), .IN3(\key_mem[11][11] ), .IN4(n7191), .Q(n5177)
          );
   AO22X1 U4390 (.IN1(n7183), .IN2(n2875), .IN3(\key_mem[12][11] ), .IN4(n7185), .Q(n5178)
          );
   AO22X1 U4391 (.IN1(n7182), .IN2(n2875), .IN3(\key_mem[13][11] ), .IN4(n7170), .Q(n5179)
          );
   AO22X1 U4392 (.IN1(n6992), .IN2(n2875), .IN3(\key_mem[14][11] ), .IN4(n7151), .Q(n5180)
          );
   AO221X1 U4393 (.IN1(n7135), .IN2(n2876), .IN3(key[139]), .IN4(n7294), .IN5(n2877), .Q(
          n2875));
   AO222X1 U4394 (.IN1(n7109), .IN2(n2878), .IN3(key[11]), .IN4(n7080), .IN5(n7047), .IN6(
          n2879), .Q(n2877));
   AO22X1 U4395 (.IN1(n7295), .IN2(n2880), .IN3(\key_mem[0][10] ), .IN4(n6928), .Q(n5181)
          );
   AO22X1 U4396 (.IN1(n6927), .IN2(n2880), .IN3(\key_mem[1][10] ), .IN4(n6825), .Q(n5182)
          );
   AO22X1 U4397 (.IN1(n6856), .IN2(n2880), .IN3(\key_mem[2][10] ), .IN4(n6849), .Q(n5183)
          );
   AO22X1 U4398 (.IN1(n6870), .IN2(n2880), .IN3(\key_mem[3][10] ), .IN4(n6863), .Q(n5184)
          );
   AO22X1 U4399 (.IN1(n6889), .IN2(n2880), .IN3(\key_mem[4][10] ), .IN4(n6890), .Q(n5185)
          );
   AO22X1 U4400 (.IN1(n7020), .IN2(n2880), .IN3(\key_mem[5][10] ), .IN4(n7270), .Q(n5186)
          );
   AO22X1 U4401 (.IN1(n6969), .IN2(n2880), .IN3(\key_mem[6][10] ), .IN4(n7252), .Q(n5187)
          );
   AO22X1 U4402 (.IN1(n7244), .IN2(n2880), .IN3(\key_mem[7][10] ), .IN4(n7242), .Q(n5188)
          );
   AO22X1 U4403 (.IN1(n6749), .IN2(n2880), .IN3(\key_mem[8][10] ), .IN4(n6721), .Q(n5189)
          );
   AO22X1 U4404 (.IN1(n7009), .IN2(n2880), .IN3(\key_mem[9][10] ), .IN4(n7213), .Q(n5190)
          );
   AO22X1 U4405 (.IN1(n6796), .IN2(n2880), .IN3(\key_mem[10][10] ), .IN4(n6768), .Q(n5191)
          );
   AO22X1 U4406 (.IN1(n7004), .IN2(n2880), .IN3(\key_mem[11][10] ), .IN4(n7189), .Q(n5192)
          );
   AO22X1 U4407 (.IN1(n7186), .IN2(n2880), .IN3(\key_mem[12][10] ), .IN4(n6983), .Q(n5193)
          );
   AO22X1 U4408 (.IN1(n6999), .IN2(n2880), .IN3(\key_mem[13][10] ), .IN4(n7168), .Q(n5194)
          );
   AO22X1 U4409 (.IN1(n7161), .IN2(n2880), .IN3(\key_mem[14][10] ), .IN4(n7150), .Q(n5195)
          );
   AO222X1 U4411 (.IN1(n7109), .IN2(n2883), .IN3(key[10]), .IN4(n7080), .IN5(n7047), .IN6(
          n2884), .Q(n2882));
   AO22X1 U4412 (.IN1(n7304), .IN2(n2885), .IN3(\key_mem[0][9] ), .IN4(n6928), .Q(n5196)
          );
   AO22X1 U4413 (.IN1(n6811), .IN2(n2885), .IN3(\key_mem[1][9] ), .IN4(n6815), .Q(n5197)
          );
   AO22X1 U4414 (.IN1(n6988), .IN2(n2885), .IN3(\key_mem[2][9] ), .IN4(n6850), .Q(n5198)
          );
   AO22X1 U4415 (.IN1(n6870), .IN2(n2885), .IN3(\key_mem[3][9] ), .IN4(n6861), .Q(n5199)
          );
   AO22X1 U4416 (.IN1(n6921), .IN2(n2885), .IN3(\key_mem[4][9] ), .IN4(n6917), .Q(n5200)
          );
   AO22X1 U4417 (.IN1(n7280), .IN2(n2885), .IN3(\key_mem[5][9] ), .IN4(n7282), .Q(n5201)
          );
   AO22X1 U4418 (.IN1(n6969), .IN2(n2885), .IN3(\key_mem[6][9] ), .IN4(n2283), .Q(n5202)
          );
   AO22X1 U4419 (.IN1(n7244), .IN2(n2885), .IN3(\key_mem[7][9] ), .IN4(n2284), .Q(n5203)
          );
   AO22X1 U4420 (.IN1(n6750), .IN2(n2885), .IN3(\key_mem[8][9] ), .IN4(n6731), .Q(n5204)
          );
   AO22X1 U4421 (.IN1(n7224), .IN2(n2885), .IN3(\key_mem[9][9] ), .IN4(n7226), .Q(n5205)
          );
   AO22X1 U4422 (.IN1(n6797), .IN2(n2885), .IN3(\key_mem[10][9] ), .IN4(n6778), .Q(n5206)
          );
   AO22X1 U4423 (.IN1(n7200), .IN2(n2885), .IN3(\key_mem[11][9] ), .IN4(n7202), .Q(n5207)
          );
   AO22X1 U4424 (.IN1(n6986), .IN2(n2885), .IN3(\key_mem[12][9] ), .IN4(n7185), .Q(n5208)
          );
   AO22X1 U4425 (.IN1(n7179), .IN2(n2885), .IN3(\key_mem[13][9] ), .IN4(n7181), .Q(n5209)
          );
   AO22X1 U4426 (.IN1(n7159), .IN2(n2885), .IN3(\key_mem[14][9] ), .IN4(n7151), .Q(n5210)
          );
   AO222X1 U4428 (.IN1(n7109), .IN2(n2888), .IN3(key[9]), .IN4(n7080), .IN5(n7047), .IN6(
          n2889), .Q(n2887));
   AO22X1 U4429 (.IN1(n7303), .IN2(n2890), .IN3(\key_mem[0][8] ), .IN4(n6928), .Q(n5211)
          );
   AO22X1 U4430 (.IN1(n6810), .IN2(n2890), .IN3(\key_mem[1][8] ), .IN4(n6814), .Q(n5212)
          );
   AO22X1 U4431 (.IN1(n6853), .IN2(n2890), .IN3(\key_mem[2][8] ), .IN4(n6845), .Q(n5213)
          );
   AO22X1 U4432 (.IN1(n6869), .IN2(n2890), .IN3(\key_mem[3][8] ), .IN4(n6865), .Q(n5214)
          );
   AO22X1 U4433 (.IN1(n6921), .IN2(n2890), .IN3(\key_mem[4][8] ), .IN4(n6890), .Q(n5215)
          );
   AO22X1 U4434 (.IN1(n7274), .IN2(n2890), .IN3(\key_mem[5][8] ), .IN4(n7270), .Q(n5216)
          );
   AO22X1 U4435 (.IN1(n6969), .IN2(n2890), .IN3(\key_mem[6][8] ), .IN4(n7259), .Q(n5217)
          );
   AO22X1 U4436 (.IN1(n7249), .IN2(n2890), .IN3(\key_mem[7][8] ), .IN4(n7241), .Q(n5218)
          );
   AO22X1 U4437 (.IN1(n6758), .IN2(n2890), .IN3(\key_mem[8][8] ), .IN4(n6741), .Q(n5219)
          );
   AO22X1 U4438 (.IN1(n7218), .IN2(n2890), .IN3(\key_mem[9][8] ), .IN4(n7214), .Q(n5220)
          );
   AO22X1 U4439 (.IN1(n6805), .IN2(n2890), .IN3(\key_mem[10][8] ), .IN4(n6788), .Q(n5221)
          );
   AO22X1 U4440 (.IN1(n7194), .IN2(n2890), .IN3(\key_mem[11][8] ), .IN4(n7190), .Q(n5222)
          );
   AO22X1 U4441 (.IN1(n6829), .IN2(n2890), .IN3(\key_mem[12][8] ), .IN4(n2289), .Q(n5223)
          );
   AO22X1 U4442 (.IN1(n7173), .IN2(n2890), .IN3(\key_mem[13][8] ), .IN4(n7169), .Q(n5224)
          );
   AO22X1 U4443 (.IN1(n7158), .IN2(n2890), .IN3(\key_mem[14][8] ), .IN4(n7148), .Q(n5225)
          );
   AO221X1 U4444 (.IN1(n7135), .IN2(n2891), .IN3(key[136]), .IN4(n7309), .IN5(n2892), .Q(
          n2890));
   AO222X1 U4445 (.IN1(n7109), .IN2(n2893), .IN3(key[8]), .IN4(n7080), .IN5(n7047), .IN6(
          n2894), .Q(n2892));
   AO22X1 U4446 (.IN1(n7297), .IN2(n2895), .IN3(\key_mem[0][7] ), .IN4(n6928), .Q(n5226)
          );
   AO22X1 U4447 (.IN1(n6811), .IN2(n2895), .IN3(\key_mem[1][7] ), .IN4(n6820), .Q(n5227)
          );
   AO22X1 U4448 (.IN1(n6856), .IN2(n2895), .IN3(\key_mem[2][7] ), .IN4(n6847), .Q(n5228)
          );
   AO22X1 U4449 (.IN1(n6874), .IN2(n2895), .IN3(\key_mem[3][7] ), .IN4(n6864), .Q(n5229)
          );
   AO22X1 U4450 (.IN1(n6888), .IN2(n2895), .IN3(\key_mem[4][7] ), .IN4(n6919), .Q(n5230)
          );
   AO22X1 U4451 (.IN1(n7276), .IN2(n2895), .IN3(\key_mem[5][7] ), .IN4(n7270), .Q(n5231)
          );
   AO22X1 U4452 (.IN1(n7261), .IN2(n2895), .IN3(\key_mem[6][7] ), .IN4(n7251), .Q(n5232)
          );
   AO22X1 U4453 (.IN1(n7245), .IN2(n2895), .IN3(\key_mem[7][7] ), .IN4(n2284), .Q(n5233)
          );
   AO22X1 U4454 (.IN1(n6748), .IN2(n2895), .IN3(\key_mem[8][7] ), .IN4(n6733), .Q(n5234)
          );
   AO22X1 U4455 (.IN1(n7220), .IN2(n2895), .IN3(\key_mem[9][7] ), .IN4(n7213), .Q(n5235)
          );
   AO22X1 U4456 (.IN1(n6795), .IN2(n2895), .IN3(\key_mem[10][7] ), .IN4(n6780), .Q(n5236)
          );
   AO22X1 U4457 (.IN1(n7196), .IN2(n2895), .IN3(\key_mem[11][7] ), .IN4(n7189), .Q(n5237)
          );
   AO22X1 U4458 (.IN1(n6832), .IN2(n2895), .IN3(\key_mem[12][7] ), .IN4(n6983), .Q(n5238)
          );
   AO22X1 U4459 (.IN1(n7175), .IN2(n2895), .IN3(\key_mem[13][7] ), .IN4(n7168), .Q(n5239)
          );
   AO22X1 U4460 (.IN1(n7161), .IN2(n2895), .IN3(\key_mem[14][7] ), .IN4(n7149), .Q(n5240)
          );
   AO221X1 U4461 (.IN1(n7136), .IN2(n2896), .IN3(key[135]), .IN4(n7305), .IN5(n2897), .Q(
          n2895));
   AO222X1 U4462 (.IN1(n7109), .IN2(n2898), .IN3(key[7]), .IN4(n7081), .IN5(n7048), .IN6(
          n2899), .Q(n2897));
   AO22X1 U4463 (.IN1(n7296), .IN2(n2900), .IN3(\key_mem[0][6] ), .IN4(n6928), .Q(n5241)
          );
   AO22X1 U4464 (.IN1(n6808), .IN2(n2900), .IN3(\key_mem[1][6] ), .IN4(n6818), .Q(n5242)
          );
   AO22X1 U4465 (.IN1(n6855), .IN2(n2900), .IN3(\key_mem[2][6] ), .IN4(n6842), .Q(n5243)
          );
   AO22X1 U4466 (.IN1(n6875), .IN2(n2900), .IN3(\key_mem[3][6] ), .IN4(n6867), .Q(n5244)
          );
   AO22X1 U4467 (.IN1(n6916), .IN2(n2900), .IN3(\key_mem[4][6] ), .IN4(n6918), .Q(n5245)
          );
   AO22X1 U4468 (.IN1(n7277), .IN2(n2900), .IN3(\key_mem[5][6] ), .IN4(n7267), .Q(n5246)
          );
   AO22X1 U4469 (.IN1(n7260), .IN2(n2900), .IN3(\key_mem[6][6] ), .IN4(n7257), .Q(n5247)
          );
   AO22X1 U4470 (.IN1(n7245), .IN2(n2900), .IN3(\key_mem[7][6] ), .IN4(n7012), .Q(n5248)
          );
   AO22X1 U4471 (.IN1(n6749), .IN2(n2900), .IN3(\key_mem[8][6] ), .IN4(n6727), .Q(n5249)
          );
   AO22X1 U4472 (.IN1(n7221), .IN2(n2900), .IN3(\key_mem[9][6] ), .IN4(n7211), .Q(n5250)
          );
   AO22X1 U4473 (.IN1(n6796), .IN2(n2900), .IN3(\key_mem[10][6] ), .IN4(n6774), .Q(n5251)
          );
   AO22X1 U4474 (.IN1(n7197), .IN2(n2900), .IN3(\key_mem[11][6] ), .IN4(n7187), .Q(n5252)
          );
   AO22X1 U4475 (.IN1(n6840), .IN2(n2900), .IN3(\key_mem[12][6] ), .IN4(n7185), .Q(n5253)
          );
   AO22X1 U4476 (.IN1(n7176), .IN2(n2900), .IN3(\key_mem[13][6] ), .IN4(n7166), .Q(n5254)
          );
   AO22X1 U4477 (.IN1(n7160), .IN2(n2900), .IN3(\key_mem[14][6] ), .IN4(n7156), .Q(n5255)
          );
   AO222X1 U4479 (.IN1(n7109), .IN2(n2903), .IN3(key[6]), .IN4(n7081), .IN5(n7048), .IN6(
          n2904), .Q(n2902));
   AO22X1 U4480 (.IN1(n7295), .IN2(n2905), .IN3(\key_mem[0][5] ), .IN4(n6928), .Q(n5256)
          );
   AO22X1 U4481 (.IN1(n6809), .IN2(n2905), .IN3(\key_mem[1][5] ), .IN4(n6821), .Q(n5257)
          );
   AO22X1 U4482 (.IN1(n6988), .IN2(n2905), .IN3(\key_mem[2][5] ), .IN4(n6842), .Q(n5258)
          );
   AO22X1 U4483 (.IN1(n6807), .IN2(n2905), .IN3(\key_mem[3][5] ), .IN4(n6862), .Q(n5259)
          );
   AO22X1 U4484 (.IN1(n7286), .IN2(n2905), .IN3(\key_mem[4][5] ), .IN4(n7284), .Q(n5260)
          );
   AO22X1 U4485 (.IN1(n7279), .IN2(n2905), .IN3(\key_mem[5][5] ), .IN4(n7268), .Q(n5261)
          );
   AO22X1 U4486 (.IN1(n7265), .IN2(n2905), .IN3(\key_mem[6][5] ), .IN4(n7254), .Q(n5262)
          );
   AO22X1 U4487 (.IN1(n7246), .IN2(n2905), .IN3(\key_mem[7][5] ), .IN4(n7243), .Q(n5263)
          );
   AO22X1 U4488 (.IN1(n6754), .IN2(n2905), .IN3(\key_mem[8][5] ), .IN4(n6715), .Q(n5264)
          );
   AO22X1 U4489 (.IN1(n7223), .IN2(n2905), .IN3(\key_mem[9][5] ), .IN4(n7212), .Q(n5265)
          );
   AO22X1 U4490 (.IN1(n6801), .IN2(n2905), .IN3(\key_mem[10][5] ), .IN4(n6762), .Q(n5266)
          );
   AO22X1 U4491 (.IN1(n7199), .IN2(n2905), .IN3(\key_mem[11][5] ), .IN4(n7188), .Q(n5267)
          );
   AO22X1 U4492 (.IN1(n6831), .IN2(n2905), .IN3(\key_mem[12][5] ), .IN4(n7000), .Q(n5268)
          );
   AO22X1 U4493 (.IN1(n7178), .IN2(n2905), .IN3(\key_mem[13][5] ), .IN4(n7167), .Q(n5269)
          );
   AO22X1 U4494 (.IN1(n7164), .IN2(n2905), .IN3(\key_mem[14][5] ), .IN4(n7157), .Q(n5270)
          );
   AO221X1 U4495 (.IN1(n7136), .IN2(n2906), .IN3(key[133]), .IN4(n7309), .IN5(n2907), .Q(
          n2905));
   AO222X1 U4496 (.IN1(n7109), .IN2(n2908), .IN3(key[5]), .IN4(n7081), .IN5(n7048), .IN6(
          n2909), .Q(n2907));
   AO22X1 U4497 (.IN1(n7304), .IN2(n2910), .IN3(\key_mem[0][4] ), .IN4(n6928), .Q(n5271)
          );
   AO22X1 U4498 (.IN1(n6810), .IN2(n2910), .IN3(\key_mem[1][4] ), .IN4(n6817), .Q(n5272)
          );
   AO22X1 U4499 (.IN1(n6856), .IN2(n2910), .IN3(\key_mem[2][4] ), .IN4(n6850), .Q(n5273)
          );
   AO22X1 U4500 (.IN1(n6872), .IN2(n2910), .IN3(\key_mem[3][4] ), .IN4(n6865), .Q(n5274)
          );
   AO22X1 U4501 (.IN1(n6888), .IN2(n2910), .IN3(\key_mem[4][4] ), .IN4(n7021), .Q(n5275)
          );
   AO22X1 U4502 (.IN1(n6974), .IN2(n2910), .IN3(\key_mem[5][4] ), .IN4(n7271), .Q(n5276)
          );
   AO22X1 U4503 (.IN1(n6970), .IN2(n2910), .IN3(\key_mem[6][4] ), .IN4(n7255), .Q(n5277)
          );
   AO22X1 U4504 (.IN1(n7247), .IN2(n2910), .IN3(\key_mem[7][4] ), .IN4(n7235), .Q(n5278)
          );
   AO22X1 U4505 (.IN1(n6755), .IN2(n2910), .IN3(\key_mem[8][4] ), .IN4(n6739), .Q(n5279)
          );
   AO22X1 U4506 (.IN1(n6976), .IN2(n2910), .IN3(\key_mem[9][4] ), .IN4(n7215), .Q(n5280)
          );
   AO22X1 U4507 (.IN1(n6802), .IN2(n2910), .IN3(\key_mem[10][4] ), .IN4(n6786), .Q(n5281)
          );
   AO22X1 U4508 (.IN1(n6978), .IN2(n2910), .IN3(\key_mem[11][4] ), .IN4(n7191), .Q(n5282)
          );
   AO22X1 U4509 (.IN1(n6827), .IN2(n2910), .IN3(\key_mem[12][4] ), .IN4(n6985), .Q(n5283)
          );
   AO22X1 U4510 (.IN1(n6980), .IN2(n2910), .IN3(\key_mem[13][4] ), .IN4(n7170), .Q(n5284)
          );
   AO22X1 U4511 (.IN1(n6972), .IN2(n2910), .IN3(\key_mem[14][4] ), .IN4(n6994), .Q(n5285)
          );
   AO222X1 U4513 (.IN1(n7108), .IN2(n2913), .IN3(key[4]), .IN4(n7081), .IN5(n7048), .IN6(
          n2914), .Q(n2912));
   AO22X1 U4514 (.IN1(n7308), .IN2(n2915), .IN3(\key_mem[0][3] ), .IN4(n6928), .Q(n5286)
          );
   AO22X1 U4515 (.IN1(n6811), .IN2(n2915), .IN3(\key_mem[1][3] ), .IN4(n6814), .Q(n5287)
          );
   AO22X1 U4516 (.IN1(n6856), .IN2(n2915), .IN3(\key_mem[2][3] ), .IN4(n6849), .Q(n5288)
          );
   AO22X1 U4517 (.IN1(n6807), .IN2(n2915), .IN3(\key_mem[3][3] ), .IN4(n6868), .Q(n5289)
          );
   AO22X1 U4518 (.IN1(n7287), .IN2(n2915), .IN3(\key_mem[4][3] ), .IN4(n6915), .Q(n5290)
          );
   AO22X1 U4519 (.IN1(n7283), .IN2(n2915), .IN3(\key_mem[5][3] ), .IN4(n7267), .Q(n5291)
          );
   AO22X1 U4520 (.IN1(n6969), .IN2(n2915), .IN3(\key_mem[6][3] ), .IN4(n7252), .Q(n5292)
          );
   AO22X1 U4521 (.IN1(n7248), .IN2(n2915), .IN3(\key_mem[7][3] ), .IN4(n7236), .Q(n5293)
          );
   AO22X1 U4522 (.IN1(n6751), .IN2(n2915), .IN3(\key_mem[8][3] ), .IN4(n6731), .Q(n5294)
          );
   AO22X1 U4523 (.IN1(n7227), .IN2(n2915), .IN3(\key_mem[9][3] ), .IN4(n7211), .Q(n5295)
          );
   AO22X1 U4524 (.IN1(n6798), .IN2(n2915), .IN3(\key_mem[10][3] ), .IN4(n6778), .Q(n5296)
          );
   AO22X1 U4525 (.IN1(n7203), .IN2(n2915), .IN3(\key_mem[11][3] ), .IN4(n7187), .Q(n5297)
          );
   AO22X1 U4526 (.IN1(n7183), .IN2(n2915), .IN3(\key_mem[12][3] ), .IN4(n7185), .Q(n5298)
          );
   AO22X1 U4527 (.IN1(n7182), .IN2(n2915), .IN3(\key_mem[13][3] ), .IN4(n7166), .Q(n5299)
          );
   AO22X1 U4528 (.IN1(n6971), .IN2(n2915), .IN3(\key_mem[14][3] ), .IN4(n7151), .Q(n5300)
          );
   AO221X1 U4529 (.IN1(n7136), .IN2(n2916), .IN3(key[131]), .IN4(n7290), .IN5(n2917), .Q(
          n2915));
   AO222X1 U4530 (.IN1(n7108), .IN2(n2918), .IN3(key[3]), .IN4(n7081), .IN5(n7048), .IN6(
          n2919), .Q(n2917));
   AO22X1 U4531 (.IN1(n7295), .IN2(n2920), .IN3(\key_mem[0][2] ), .IN4(n6928), .Q(n5301)
          );
   AO22X1 U4532 (.IN1(n6926), .IN2(n2920), .IN3(\key_mem[1][2] ), .IN4(n6815), .Q(n5302)
          );
   AO22X1 U4533 (.IN1(n6853), .IN2(n2920), .IN3(\key_mem[2][2] ), .IN4(n6847), .Q(n5303)
          );
   AO22X1 U4534 (.IN1(n6874), .IN2(n2920), .IN3(\key_mem[3][2] ), .IN4(n6865), .Q(n5304)
          );
   AO22X1 U4535 (.IN1(n7287), .IN2(n2920), .IN3(\key_mem[4][2] ), .IN4(n7285), .Q(n5305)
          );
   AO22X1 U4536 (.IN1(n7283), .IN2(n2920), .IN3(\key_mem[5][2] ), .IN4(n7271), .Q(n5306)
          );
   AO22X1 U4537 (.IN1(n7261), .IN2(n2920), .IN3(\key_mem[6][2] ), .IN4(n7253), .Q(n5307)
          );
   AO22X1 U4538 (.IN1(n7250), .IN2(n2920), .IN3(\key_mem[7][2] ), .IN4(n7237), .Q(n5308)
          );
   AO22X1 U4539 (.IN1(n6752), .IN2(n2920), .IN3(\key_mem[8][2] ), .IN4(n6725), .Q(n5309)
          );
   AO22X1 U4540 (.IN1(n7227), .IN2(n2920), .IN3(\key_mem[9][2] ), .IN4(n7215), .Q(n5310)
          );
   AO22X1 U4541 (.IN1(n6799), .IN2(n2920), .IN3(\key_mem[10][2] ), .IN4(n6772), .Q(n5311)
          );
   AO22X1 U4542 (.IN1(n7203), .IN2(n2920), .IN3(\key_mem[11][2] ), .IN4(n7191), .Q(n5312)
          );
   AO22X1 U4543 (.IN1(n6829), .IN2(n2920), .IN3(\key_mem[12][2] ), .IN4(n6984), .Q(n5313)
          );
   AO22X1 U4544 (.IN1(n7182), .IN2(n2920), .IN3(\key_mem[13][2] ), .IN4(n7170), .Q(n5314)
          );
   AO22X1 U4545 (.IN1(n6971), .IN2(n2920), .IN3(\key_mem[14][2] ), .IN4(n7152), .Q(n5315)
          );
   AO221X1 U4546 (.IN1(n7136), .IN2(n2921), .IN3(key[130]), .IN4(n7294), .IN5(n2922), .Q(
          n2920));
   AO222X1 U4547 (.IN1(n7108), .IN2(n2923), .IN3(key[2]), .IN4(n7081), .IN5(n7048), .IN6(
          n2924), .Q(n2922));
   AO22X1 U4548 (.IN1(n7311), .IN2(n2925), .IN3(\key_mem[0][1] ), .IN4(n6928), .Q(n5316)
          );
   AO22X1 U4549 (.IN1(n6811), .IN2(n2925), .IN3(\key_mem[1][1] ), .IN4(n6816), .Q(n5317)
          );
   AO22X1 U4550 (.IN1(n6854), .IN2(n2925), .IN3(\key_mem[2][1] ), .IN4(n6849), .Q(n5318)
          );
   AO22X1 U4551 (.IN1(n6875), .IN2(n2925), .IN3(\key_mem[3][1] ), .IN4(n6865), .Q(n5319)
          );
   AO22X1 U4552 (.IN1(n7286), .IN2(n2925), .IN3(\key_mem[4][1] ), .IN4(n6919), .Q(n5320)
          );
   AO22X1 U4553 (.IN1(n7019), .IN2(n2925), .IN3(\key_mem[5][1] ), .IN4(n2282), .Q(n5321)
          );
   AO22X1 U4554 (.IN1(n7263), .IN2(n2925), .IN3(\key_mem[6][1] ), .IN4(n7252), .Q(n5322)
          );
   AO22X1 U4555 (.IN1(n7245), .IN2(n2925), .IN3(\key_mem[7][1] ), .IN4(n7238), .Q(n5323)
          );
   AO22X1 U4556 (.IN1(n6754), .IN2(n2925), .IN3(\key_mem[8][1] ), .IN4(n6714), .Q(n5324)
          );
   AO22X1 U4557 (.IN1(n7008), .IN2(n2925), .IN3(\key_mem[9][1] ), .IN4(n2286), .Q(n5325)
          );
   AO22X1 U4558 (.IN1(n6801), .IN2(n2925), .IN3(\key_mem[10][1] ), .IN4(n6761), .Q(n5326)
          );
   AO22X1 U4559 (.IN1(n7003), .IN2(n2925), .IN3(\key_mem[11][1] ), .IN4(n2288), .Q(n5327)
          );
   AO22X1 U4560 (.IN1(n6829), .IN2(n2925), .IN3(\key_mem[12][1] ), .IN4(n6983), .Q(n5328)
          );
   AO22X1 U4561 (.IN1(n6998), .IN2(n2925), .IN3(\key_mem[13][1] ), .IN4(n2290), .Q(n5329)
          );
   AO22X1 U4562 (.IN1(n6992), .IN2(n2925), .IN3(\key_mem[14][1] ), .IN4(n7153), .Q(n5330)
          );
   AO222X1 U4564 (.IN1(n7108), .IN2(n2928), .IN3(key[1]), .IN4(n7081), .IN5(n7048), .IN6(
          n2929), .Q(n2927));
   AO22X1 U4565 (.IN1(n7290), .IN2(n2930), .IN3(\key_mem[0][0] ), .IN4(n6928), .Q(n5331)
          );
   AO22X1 U4566 (.IN1(n6927), .IN2(n2930), .IN3(\key_mem[1][0] ), .IN4(n6816), .Q(n5332)
          );
   AO22X1 U4567 (.IN1(n6855), .IN2(n2930), .IN3(\key_mem[2][0] ), .IN4(n6851), .Q(n5333)
          );
   AO22X1 U4568 (.IN1(n6873), .IN2(n2930), .IN3(\key_mem[3][0] ), .IN4(n6866), .Q(n5334)
          );
   NOR3X0 U4569 (.IN1(round_ctr_reg[2]), .IN2(round_ctr_reg[3]), .IN3(n2213), .QN(n2932)
          );
   AO22X1 U4570 (.IN1(n7286), .IN2(n2930), .IN3(\key_mem[4][0] ), .IN4(n7021), .Q(n5335)
          );
   AO22X1 U4572 (.IN1(n7278), .IN2(n2930), .IN3(\key_mem[5][0] ), .IN4(n7282), .Q(n5336)
          );
   AO22X1 U4574 (.IN1(n7262), .IN2(n2930), .IN3(\key_mem[6][0] ), .IN4(n2283), .Q(n5337)
          );
   AO22X1 U4575 (.IN1(n7245), .IN2(n2930), .IN3(\key_mem[7][0] ), .IN4(n7239), .Q(n5338)
          );
   AO22X1 U4576 (.IN1(n6755), .IN2(n2930), .IN3(\key_mem[8][0] ), .IN4(n6720), .Q(n5339)
          );
   AO22X1 U4578 (.IN1(n7222), .IN2(n2930), .IN3(\key_mem[9][0] ), .IN4(n7226), .Q(n5340)
          );
   AO22X1 U4580 (.IN1(n6802), .IN2(n2930), .IN3(\key_mem[10][0] ), .IN4(n6767), .Q(n5341)
          );
   AO22X1 U4582 (.IN1(n7198), .IN2(n2930), .IN3(\key_mem[11][0] ), .IN4(n7202), .Q(n5342)
          );
   AO22X1 U4584 (.IN1(n6832), .IN2(n2930), .IN3(\key_mem[12][0] ), .IN4(n6839), .Q(n5343)
          );
   AO22X1 U4586 (.IN1(n7177), .IN2(n2930), .IN3(\key_mem[13][0] ), .IN4(n7181), .Q(n5344)
          );
   AO22X1 U4589 (.IN1(n7159), .IN2(n2930), .IN3(\key_mem[14][0] ), .IN4(n7150), .Q(n5345)
          );
   AO221X1 U4590 (.IN1(n7136), .IN2(n2937), .IN3(key[128]), .IN4(n2276), .IN5(n2938), .Q(
          n2930));
   AO222X1 U4591 (.IN1(n7108), .IN2(n2939), .IN3(key[0]), .IN4(n7081), .IN5(n7048), .IN6(
          n2940), .Q(n2938));
   AOI222X1 U4593 (.IN1(n2299), .IN2(n7048), .IN3(n2293), .IN4(n7136), .IN5(n2296), .IN6(
          n7108), .QN(n2943));
   XNOR2X1 U4594 (.IN1(prev_key0_reg[127]), .IN2(n7590), .Q(n2296));
   XNOR2X1 U4595 (.IN1(prev_key0_reg[127]), .IN2(n7598), .Q(n2293));
   XNOR2X1 U4596 (.IN1(prev_key1_reg[127]), .IN2(n7590), .Q(n2299));
   AOI222X1 U4597 (.IN1(prev_key1_reg[127]), .IN2(n6951), .IN3(n7081), .IN4(key[127]), .
          IN5(key[255]), .IN6(n6704), .QN(n2942));
   AOI222X1 U4598 (.IN1(n2304), .IN2(n7048), .IN3(n2301), .IN4(n7136), .IN5(n2303), .IN6(
          n7108), .QN(n2947));
   XNOR2X1 U4599 (.IN1(prev_key0_reg[126]), .IN2(n2948), .Q(n2303));
   XNOR2X1 U4600 (.IN1(prev_key0_reg[126]), .IN2(n7597), .Q(n2301));
   XNOR2X1 U4601 (.IN1(prev_key1_reg[126]), .IN2(n2948), .Q(n2304));
   AOI222X1 U4602 (.IN1(prev_key1_reg[126]), .IN2(n6949), .IN3(n7081), .IN4(key[126]), .
          IN5(key[254]), .IN6(n6703), .QN(n2946));
   AOI222X1 U4603 (.IN1(n2309), .IN2(n7048), .IN3(n2306), .IN4(n7136), .IN5(n2308), .IN6(
          n7108), .QN(n2950));
   XNOR2X1 U4604 (.IN1(prev_key0_reg[125]), .IN2(n2951), .Q(n2308));
   XNOR2X1 U4605 (.IN1(prev_key0_reg[125]), .IN2(n7596), .Q(n2306));
   XNOR2X1 U4606 (.IN1(prev_key1_reg[125]), .IN2(n2951), .Q(n2309));
   AOI222X1 U4607 (.IN1(prev_key1_reg[125]), .IN2(n6945), .IN3(n7081), .IN4(key[125]), .
          IN5(key[253]), .IN6(n6710), .QN(n2949));
   AOI222X1 U4608 (.IN1(n2314), .IN2(n7048), .IN3(n2311), .IN4(n7136), .IN5(n2313), .IN6(
          n7108), .QN(n2953));
   XNOR2X1 U4609 (.IN1(prev_key0_reg[124]), .IN2(n2954), .Q(n2313));
   XNOR2X1 U4610 (.IN1(prev_key0_reg[124]), .IN2(n7595), .Q(n2311));
   XNOR2X1 U4611 (.IN1(prev_key1_reg[124]), .IN2(n2954), .Q(n2314));
   AOI222X1 U4612 (.IN1(prev_key1_reg[124]), .IN2(n6947), .IN3(n7081), .IN4(key[124]), .
          IN5(key[252]), .IN6(n6709), .QN(n2952));
   AOI222X1 U4613 (.IN1(n2319), .IN2(n7048), .IN3(n2316), .IN4(n7136), .IN5(n2318), .IN6(
          n7108), .QN(n2956));
   XNOR2X1 U4614 (.IN1(prev_key0_reg[123]), .IN2(n2957), .Q(n2318));
   XNOR2X1 U4615 (.IN1(prev_key0_reg[123]), .IN2(n7594), .Q(n2316));
   XNOR2X1 U4616 (.IN1(prev_key1_reg[123]), .IN2(n2957), .Q(n2319));
   AOI222X1 U4617 (.IN1(prev_key1_reg[123]), .IN2(n6952), .IN3(n7081), .IN4(key[123]), .
          IN5(key[251]), .IN6(n6708), .QN(n2955));
   AOI222X1 U4618 (.IN1(n2324), .IN2(n7048), .IN3(n2321), .IN4(n7137), .IN5(n2323), .IN6(
          n7108), .QN(n2959));
   XNOR2X1 U4619 (.IN1(prev_key0_reg[122]), .IN2(n2960), .Q(n2323));
   XNOR2X1 U4620 (.IN1(prev_key0_reg[122]), .IN2(n7593), .Q(n2321));
   XNOR2X1 U4621 (.IN1(prev_key1_reg[122]), .IN2(n2960), .Q(n2324));
   AOI222X1 U4622 (.IN1(prev_key1_reg[122]), .IN2(n6950), .IN3(n7082), .IN4(key[122]), .
          IN5(key[250]), .IN6(n6707), .QN(n2958));
   AOI222X1 U4623 (.IN1(n2329), .IN2(n7049), .IN3(n2326), .IN4(n7137), .IN5(n2328), .IN6(
          n7108), .QN(n2962));
   XNOR2X1 U4624 (.IN1(prev_key0_reg[121]), .IN2(n2963), .Q(n2328));
   XNOR2X1 U4625 (.IN1(prev_key0_reg[121]), .IN2(n7592), .Q(n2326));
   XNOR2X1 U4626 (.IN1(prev_key1_reg[121]), .IN2(n2963), .Q(n2329));
   AOI222X1 U4627 (.IN1(prev_key1_reg[121]), .IN2(n6955), .IN3(n7082), .IN4(key[121]), .
          IN5(key[249]), .IN6(n6706), .QN(n2961));
   AOI222X1 U4628 (.IN1(n2334), .IN2(n7049), .IN3(n2331), .IN4(n7137), .IN5(n2333), .IN6(
          n7108), .QN(n2965));
   XNOR2X1 U4629 (.IN1(prev_key0_reg[120]), .IN2(n2966), .Q(n2333));
   XNOR2X1 U4630 (.IN1(prev_key0_reg[120]), .IN2(n7591), .Q(n2331));
   XNOR2X1 U4631 (.IN1(prev_key1_reg[120]), .IN2(n2966), .Q(n2334));
   AOI222X1 U4632 (.IN1(prev_key1_reg[120]), .IN2(n6950), .IN3(n7082), .IN4(key[120]), .
          IN5(key[248]), .IN6(n6705), .QN(n2964));
   AOI222X1 U4633 (.IN1(n2339), .IN2(n7049), .IN3(n2336), .IN4(n7137), .IN5(n2338), .IN6(
          n7107), .QN(n2968));
   XNOR2X1 U4634 (.IN1(prev_key0_reg[119]), .IN2(n7611), .Q(n2338));
   XNOR2X1 U4635 (.IN1(new_sboxw[23]), .IN2(n2223), .Q(n2336));
   XNOR2X1 U4636 (.IN1(prev_key1_reg[119]), .IN2(n7611), .Q(n2339));
   AOI222X1 U4637 (.IN1(prev_key1_reg[119]), .IN2(n6951), .IN3(n7082), .IN4(key[119]), .
          IN5(key[247]), .IN6(n6704), .QN(n2967));
   AOI222X1 U4638 (.IN1(n2344), .IN2(n7049), .IN3(n2341), .IN4(n7137), .IN5(n2343), .IN6(
          n7107), .QN(n2970));
   XNOR2X1 U4639 (.IN1(prev_key0_reg[118]), .IN2(n6699), .Q(n2343));
   XNOR2X1 U4641 (.IN1(prev_key1_reg[118]), .IN2(n6699), .Q(n2344));
   AOI222X1 U4642 (.IN1(prev_key1_reg[118]), .IN2(n6952), .IN3(n7082), .IN4(key[118]), .
          IN5(key[246]), .IN6(n6703), .QN(n2969));
   AOI222X1 U4643 (.IN1(n2349), .IN2(n7049), .IN3(n2346), .IN4(n7137), .IN5(n2348), .IN6(
          n7107), .QN(n2972));
   XNOR2X1 U4644 (.IN1(prev_key0_reg[117]), .IN2(n7609), .Q(n2348));
   XNOR2X1 U4645 (.IN1(new_sboxw[21]), .IN2(n2225), .Q(n2346));
   XNOR2X1 U4646 (.IN1(prev_key1_reg[117]), .IN2(n7609), .Q(n2349));
   AOI222X1 U4647 (.IN1(prev_key1_reg[117]), .IN2(n6953), .IN3(n7082), .IN4(key[117]), .
          IN5(key[245]), .IN6(n6711), .QN(n2971));
   AOI222X1 U4648 (.IN1(n2354), .IN2(n7049), .IN3(n2351), .IN4(n7137), .IN5(n2353), .IN6(
          n7107), .QN(n2974));
   XNOR2X1 U4649 (.IN1(prev_key0_reg[116]), .IN2(n7608), .Q(n2353));
   XNOR2X1 U4650 (.IN1(new_sboxw[20]), .IN2(n2226), .Q(n2351));
   XNOR2X1 U4651 (.IN1(prev_key1_reg[116]), .IN2(n7608), .Q(n2354));
   AOI222X1 U4652 (.IN1(prev_key1_reg[116]), .IN2(n6954), .IN3(n7082), .IN4(key[116]), .
          IN5(key[244]), .IN6(n2945), .QN(n2973));
   AOI222X1 U4653 (.IN1(n2359), .IN2(n7049), .IN3(n2356), .IN4(n7137), .IN5(n2358), .IN6(
          n7107), .QN(n2976));
   XNOR2X1 U4654 (.IN1(prev_key0_reg[115]), .IN2(n7607), .Q(n2358));
   XNOR2X1 U4655 (.IN1(new_sboxw[19]), .IN2(n2227), .Q(n2356));
   XNOR2X1 U4656 (.IN1(prev_key1_reg[115]), .IN2(n7607), .Q(n2359));
   AOI222X1 U4657 (.IN1(prev_key1_reg[115]), .IN2(n6946), .IN3(n7082), .IN4(key[115]), .
          IN5(key[243]), .IN6(n6711), .QN(n2975));
   AOI222X1 U4658 (.IN1(n2364), .IN2(n7049), .IN3(n2361), .IN4(n7137), .IN5(n2363), .IN6(
          n7107), .QN(n2978));
   XNOR2X1 U4659 (.IN1(prev_key0_reg[114]), .IN2(n7606), .Q(n2363));
   XNOR2X1 U4660 (.IN1(new_sboxw[18]), .IN2(n2228), .Q(n2361));
   XNOR2X1 U4661 (.IN1(prev_key1_reg[114]), .IN2(n7606), .Q(n2364));
   AOI222X1 U4662 (.IN1(prev_key1_reg[114]), .IN2(n6945), .IN3(n7082), .IN4(key[114]), .
          IN5(key[242]), .IN6(n2945), .QN(n2977));
   AOI222X1 U4663 (.IN1(n2369), .IN2(n7049), .IN3(n2366), .IN4(n7137), .IN5(n2368), .IN6(
          n7107), .QN(n2980));
   XNOR2X1 U4664 (.IN1(prev_key0_reg[113]), .IN2(n7613), .Q(n2368));
   XNOR2X1 U4665 (.IN1(new_sboxw[17]), .IN2(n2229), .Q(n2366));
   XNOR2X1 U4666 (.IN1(prev_key1_reg[113]), .IN2(n7613), .Q(n2369));
   AOI222X1 U4667 (.IN1(prev_key1_reg[113]), .IN2(n6955), .IN3(n7082), .IN4(key[113]), .
          IN5(key[241]), .IN6(n6710), .QN(n2979));
   AOI222X1 U4668 (.IN1(n2374), .IN2(n7049), .IN3(n2371), .IN4(n7137), .IN5(n2373), .IN6(
          n7107), .QN(n2982));
   XNOR2X1 U4669 (.IN1(prev_key0_reg[112]), .IN2(n7612), .Q(n2373));
   XNOR2X1 U4670 (.IN1(new_sboxw[16]), .IN2(n2230), .Q(n2371));
   XNOR2X1 U4671 (.IN1(prev_key1_reg[112]), .IN2(n7612), .Q(n2374));
   AOI222X1 U4672 (.IN1(prev_key1_reg[112]), .IN2(n6952), .IN3(n7082), .IN4(key[112]), .
          IN5(key[240]), .IN6(n6709), .QN(n2981));
   AOI222X1 U4673 (.IN1(n2379), .IN2(n7049), .IN3(n2376), .IN4(n7137), .IN5(n2378), .IN6(
          n7107), .QN(n2984));
   XNOR2X1 U4674 (.IN1(prev_key0_reg[111]), .IN2(n7621), .Q(n2378));
   XNOR2X1 U4675 (.IN1(prev_key0_reg[111]), .IN2(n7611), .Q(n2376));
   XNOR2X1 U4676 (.IN1(prev_key1_reg[111]), .IN2(n7621), .Q(n2379));
   AOI222X1 U4677 (.IN1(prev_key1_reg[111]), .IN2(n6951), .IN3(n7082), .IN4(key[111]), .
          IN5(key[239]), .IN6(n6708), .QN(n2983));
   AOI222X1 U4678 (.IN1(n2384), .IN2(n7049), .IN3(n2381), .IN4(n7137), .IN5(n2383), .IN6(
          n7107), .QN(n2986));
   XNOR2X1 U4679 (.IN1(prev_key0_reg[110]), .IN2(n7620), .Q(n2383));
   XNOR2X1 U4680 (.IN1(prev_key0_reg[110]), .IN2(n6700), .Q(n2381));
   XNOR2X1 U4681 (.IN1(prev_key1_reg[110]), .IN2(n7620), .Q(n2384));
   AOI222X1 U4682 (.IN1(prev_key1_reg[110]), .IN2(n6950), .IN3(n7082), .IN4(key[110]), .
          IN5(key[238]), .IN6(n6707), .QN(n2985));
   AOI222X1 U4683 (.IN1(n2389), .IN2(n7049), .IN3(n2386), .IN4(n7138), .IN5(n2388), .IN6(
          n7107), .QN(n2988));
   XNOR2X1 U4684 (.IN1(prev_key0_reg[109]), .IN2(n7619), .Q(n2388));
   XNOR2X1 U4685 (.IN1(prev_key0_reg[109]), .IN2(n7609), .Q(n2386));
   XNOR2X1 U4686 (.IN1(prev_key1_reg[109]), .IN2(n7619), .Q(n2389));
   AOI222X1 U4687 (.IN1(prev_key1_reg[109]), .IN2(n6944), .IN3(n7082), .IN4(key[109]), .
          IN5(key[237]), .IN6(n6706), .QN(n2987));
   AOI222X1 U4688 (.IN1(n2394), .IN2(n7049), .IN3(n2391), .IN4(n7138), .IN5(n2393), .IN6(
          n7107), .QN(n2990));
   XNOR2X1 U4689 (.IN1(prev_key0_reg[108]), .IN2(n7618), .Q(n2393));
   XNOR2X1 U4690 (.IN1(prev_key0_reg[108]), .IN2(n7608), .Q(n2391));
   XNOR2X1 U4691 (.IN1(prev_key1_reg[108]), .IN2(n7618), .Q(n2394));
   AOI222X1 U4692 (.IN1(prev_key1_reg[108]), .IN2(n6952), .IN3(n7083), .IN4(key[108]), .
          IN5(key[236]), .IN6(n6705), .QN(n2989));
   AOI222X1 U4693 (.IN1(n2399), .IN2(n7049), .IN3(n2396), .IN4(n7138), .IN5(n2398), .IN6(
          n7106), .QN(n2992));
   XNOR2X1 U4694 (.IN1(prev_key0_reg[107]), .IN2(n7617), .Q(n2398));
   XNOR2X1 U4695 (.IN1(prev_key0_reg[107]), .IN2(n7607), .Q(n2396));
   XNOR2X1 U4696 (.IN1(prev_key1_reg[107]), .IN2(n7617), .Q(n2399));
   AOI222X1 U4697 (.IN1(prev_key1_reg[107]), .IN2(n6955), .IN3(n7083), .IN4(key[107]), .
          IN5(key[235]), .IN6(n6710), .QN(n2991));
   AOI222X1 U4698 (.IN1(n2404), .IN2(n7049), .IN3(n2401), .IN4(n7138), .IN5(n2403), .IN6(
          n7106), .QN(n2994));
   XNOR2X1 U4699 (.IN1(prev_key0_reg[106]), .IN2(n7616), .Q(n2403));
   XNOR2X1 U4700 (.IN1(prev_key0_reg[106]), .IN2(n7606), .Q(n2401));
   XNOR2X1 U4701 (.IN1(prev_key1_reg[106]), .IN2(n7616), .Q(n2404));
   AOI222X1 U4702 (.IN1(prev_key1_reg[106]), .IN2(n6949), .IN3(n7083), .IN4(key[106]), .
          IN5(key[234]), .IN6(n6709), .QN(n2993));
   AOI222X1 U4703 (.IN1(n2409), .IN2(n7049), .IN3(n2406), .IN4(n7138), .IN5(n2408), .IN6(
          n7106), .QN(n2996));
   XNOR2X1 U4704 (.IN1(prev_key0_reg[105]), .IN2(n7615), .Q(n2408));
   XNOR2X1 U4705 (.IN1(prev_key0_reg[105]), .IN2(n7613), .Q(n2406));
   XNOR2X1 U4706 (.IN1(prev_key1_reg[105]), .IN2(n7615), .Q(n2409));
   AOI222X1 U4707 (.IN1(prev_key1_reg[105]), .IN2(n6944), .IN3(n7083), .IN4(key[105]), .
          IN5(key[233]), .IN6(n6704), .QN(n2995));
   AOI222X1 U4708 (.IN1(n2414), .IN2(n7050), .IN3(n2411), .IN4(n7138), .IN5(n2413), .IN6(
          n7106), .QN(n2998));
   XNOR2X1 U4709 (.IN1(prev_key0_reg[104]), .IN2(n7614), .Q(n2413));
   XNOR2X1 U4710 (.IN1(prev_key0_reg[104]), .IN2(n7612), .Q(n2411));
   XNOR2X1 U4711 (.IN1(prev_key1_reg[104]), .IN2(n7614), .Q(n2414));
   AOI222X1 U4712 (.IN1(prev_key1_reg[104]), .IN2(n6945), .IN3(n7083), .IN4(key[104]), .
          IN5(key[232]), .IN6(n6703), .QN(n2997));
   AOI222X1 U4713 (.IN1(n2419), .IN2(n7050), .IN3(n2416), .IN4(n7138), .IN5(n2418), .IN6(
          n7106), .QN(n3000));
   XNOR2X1 U4714 (.IN1(prev_key0_reg[103]), .IN2(n7598), .Q(n2418));
   XNOR2X1 U4715 (.IN1(prev_key0_reg[103]), .IN2(n7621), .Q(n2416));
   XNOR2X1 U4716 (.IN1(prev_key1_reg[103]), .IN2(n7598), .Q(n2419));
   AOI222X1 U4717 (.IN1(prev_key1_reg[103]), .IN2(n6946), .IN3(n7083), .IN4(key[103]), .
          IN5(key[231]), .IN6(n6711), .QN(n2999));
   AOI222X1 U4718 (.IN1(n2424), .IN2(n7050), .IN3(n2421), .IN4(n7138), .IN5(n2423), .IN6(
          n7106), .QN(n3002));
   XNOR2X1 U4719 (.IN1(prev_key0_reg[102]), .IN2(n7597), .Q(n2423));
   XNOR2X1 U4720 (.IN1(prev_key0_reg[102]), .IN2(n7620), .Q(n2421));
   XNOR2X1 U4721 (.IN1(prev_key1_reg[102]), .IN2(n7597), .Q(n2424));
   AOI222X1 U4722 (.IN1(prev_key1_reg[102]), .IN2(n6945), .IN3(n7083), .IN4(key[102]), .
          IN5(key[230]), .IN6(n2945), .QN(n3001));
   AOI222X1 U4723 (.IN1(n2429), .IN2(n7050), .IN3(n2426), .IN4(n7138), .IN5(n2428), .IN6(
          n7106), .QN(n3004));
   XNOR2X1 U4724 (.IN1(prev_key0_reg[101]), .IN2(n7596), .Q(n2428));
   XNOR2X1 U4725 (.IN1(prev_key0_reg[101]), .IN2(n7619), .Q(n2426));
   XNOR2X1 U4726 (.IN1(prev_key1_reg[101]), .IN2(n7596), .Q(n2429));
   AOI222X1 U4727 (.IN1(prev_key1_reg[101]), .IN2(n6946), .IN3(n7083), .IN4(key[101]), .
          IN5(key[229]), .IN6(n6710), .QN(n3003));
   AOI222X1 U4728 (.IN1(n2434), .IN2(n7050), .IN3(n2431), .IN4(n7138), .IN5(n2433), .IN6(
          n7106), .QN(n3006));
   XNOR2X1 U4729 (.IN1(prev_key0_reg[100]), .IN2(n7595), .Q(n2433));
   XNOR2X1 U4730 (.IN1(prev_key0_reg[100]), .IN2(n7618), .Q(n2431));
   XNOR2X1 U4731 (.IN1(prev_key1_reg[100]), .IN2(n7595), .Q(n2434));
   AOI222X1 U4732 (.IN1(prev_key1_reg[100]), .IN2(n6947), .IN3(n7083), .IN4(key[100]), .
          IN5(key[228]), .IN6(n6709), .QN(n3005));
   AOI222X1 U4733 (.IN1(n2439), .IN2(n7050), .IN3(n2436), .IN4(n7138), .IN5(n2438), .IN6(
          n7106), .QN(n3008));
   XNOR2X1 U4734 (.IN1(prev_key0_reg[99]), .IN2(n7594), .Q(n2438));
   XNOR2X1 U4735 (.IN1(prev_key0_reg[99]), .IN2(n7617), .Q(n2436));
   XNOR2X1 U4736 (.IN1(prev_key1_reg[99]), .IN2(n7594), .Q(n2439));
   AOI222X1 U4737 (.IN1(prev_key1_reg[99]), .IN2(n6948), .IN3(n7083), .IN4(key[99]), .IN5(
          key[227]), .IN6(n6708), .QN(n3007));
   AOI222X1 U4738 (.IN1(n2444), .IN2(n7050), .IN3(n2441), .IN4(n7138), .IN5(n2443), .IN6(
          n7106), .QN(n3010));
   XNOR2X1 U4739 (.IN1(prev_key0_reg[98]), .IN2(n7593), .Q(n2443));
   XNOR2X1 U4740 (.IN1(prev_key0_reg[98]), .IN2(n7616), .Q(n2441));
   XNOR2X1 U4741 (.IN1(prev_key1_reg[98]), .IN2(n7593), .Q(n2444));
   AOI222X1 U4742 (.IN1(prev_key1_reg[98]), .IN2(n6949), .IN3(n7083), .IN4(key[98]), .IN5(
          key[226]), .IN6(n6707), .QN(n3009));
   AOI222X1 U4743 (.IN1(n2449), .IN2(n7050), .IN3(n2446), .IN4(n7138), .IN5(n2448), .IN6(
          n7106), .QN(n3012));
   XNOR2X1 U4744 (.IN1(prev_key0_reg[97]), .IN2(n7592), .Q(n2448));
   XNOR2X1 U4745 (.IN1(prev_key0_reg[97]), .IN2(n7615), .Q(n2446));
   XNOR2X1 U4746 (.IN1(prev_key1_reg[97]), .IN2(n7592), .Q(n2449));
   AOI222X1 U4747 (.IN1(prev_key1_reg[97]), .IN2(n6953), .IN3(n7083), .IN4(key[97]), .IN5(
          key[225]), .IN6(n6708), .QN(n3011));
   AOI222X1 U4748 (.IN1(n2454), .IN2(n7050), .IN3(n2451), .IN4(n7139), .IN5(n2453), .IN6(
          n7106), .QN(n3014));
   XNOR2X1 U4749 (.IN1(prev_key0_reg[96]), .IN2(n7591), .Q(n2453));
   XNOR2X1 U4750 (.IN1(prev_key0_reg[96]), .IN2(n7614), .Q(n2451));
   XNOR2X1 U4751 (.IN1(prev_key1_reg[96]), .IN2(n7591), .Q(n2454));
   AOI222X1 U4752 (.IN1(prev_key1_reg[96]), .IN2(n6950), .IN3(n7083), .IN4(key[96]), .IN5(
          key[224]), .IN6(n6707), .QN(n3013));
   AOI222X1 U4753 (.IN1(n2459), .IN2(n7050), .IN3(n2456), .IN4(n7139), .IN5(n2458), .IN6(
          n7105), .QN(n3016));
   XNOR2X1 U4754 (.IN1(n3017), .IN2(n7590), .Q(n2458));
   XNOR2X1 U4755 (.IN1(n7598), .IN2(n3017), .Q(n2456));
   XNOR2X1 U4756 (.IN1(prev_key0_reg[95]), .IN2(n2215), .Q(n3017));
   XOR3X1 U4757 (.IN1(prev_key1_reg[95]), .IN2(prev_key1_reg[127]), .IN3(n3018), .Q(n2459)
          );
   AOI222X1 U4758 (.IN1(prev_key1_reg[95]), .IN2(n6951), .IN3(n7083), .IN4(key[95]), .IN5(
          key[223]), .IN6(n6706), .QN(n3015));
   AOI222X1 U4759 (.IN1(n2464), .IN2(n7050), .IN3(n2461), .IN4(n7139), .IN5(n2463), .IN6(
          n7105), .QN(n3020));
   XNOR2X1 U4760 (.IN1(n3021), .IN2(n2948), .Q(n2463));
   XNOR2X1 U4761 (.IN1(n7597), .IN2(n3021), .Q(n2461));
   XNOR2X1 U4762 (.IN1(prev_key0_reg[94]), .IN2(n2216), .Q(n3021));
   XOR3X1 U4763 (.IN1(prev_key1_reg[94]), .IN2(prev_key1_reg[126]), .IN3(n7589), .Q(n2464)
          );
   AOI222X1 U4764 (.IN1(prev_key1_reg[94]), .IN2(n6952), .IN3(n7084), .IN4(key[94]), .IN5(
          key[222]), .IN6(n6705), .QN(n3019));
   AOI222X1 U4765 (.IN1(n2469), .IN2(n7050), .IN3(n2466), .IN4(n7139), .IN5(n2468), .IN6(
          n7105), .QN(n3023));
   XNOR2X1 U4766 (.IN1(n3024), .IN2(n2951), .Q(n2468));
   XNOR2X1 U4767 (.IN1(n7596), .IN2(n3024), .Q(n2466));
   XNOR2X1 U4768 (.IN1(prev_key0_reg[93]), .IN2(n2217), .Q(n3024));
   XOR3X1 U4769 (.IN1(prev_key1_reg[93]), .IN2(prev_key1_reg[125]), .IN3(n7588), .Q(n2469)
          );
   AOI222X1 U4770 (.IN1(prev_key1_reg[93]), .IN2(n6953), .IN3(n7084), .IN4(key[93]), .IN5(
          key[221]), .IN6(n6704), .QN(n3022));
   AOI222X1 U4771 (.IN1(n2474), .IN2(n7050), .IN3(n2471), .IN4(n7139), .IN5(n2473), .IN6(
          n7105), .QN(n3026));
   XNOR2X1 U4772 (.IN1(n3027), .IN2(n2954), .Q(n2473));
   XNOR2X1 U4773 (.IN1(n7595), .IN2(n3027), .Q(n2471));
   XNOR2X1 U4774 (.IN1(prev_key0_reg[92]), .IN2(n2218), .Q(n3027));
   XOR3X1 U4775 (.IN1(prev_key1_reg[92]), .IN2(prev_key1_reg[124]), .IN3(n7587), .Q(n2474)
          );
   AOI222X1 U4776 (.IN1(prev_key1_reg[92]), .IN2(n6954), .IN3(n7084), .IN4(key[92]), .IN5(
          key[220]), .IN6(n6703), .QN(n3025));
   AOI222X1 U4777 (.IN1(n2479), .IN2(n7050), .IN3(n2476), .IN4(n7139), .IN5(n2478), .IN6(
          n7105), .QN(n3029));
   XNOR2X1 U4778 (.IN1(n3030), .IN2(n2957), .Q(n2478));
   XNOR2X1 U4779 (.IN1(n7594), .IN2(n3030), .Q(n2476));
   XNOR2X1 U4780 (.IN1(prev_key0_reg[91]), .IN2(n2219), .Q(n3030));
   XOR3X1 U4781 (.IN1(prev_key1_reg[91]), .IN2(prev_key1_reg[123]), .IN3(n7586), .Q(n2479)
          );
   AOI222X1 U4782 (.IN1(prev_key1_reg[91]), .IN2(n6949), .IN3(n7084), .IN4(key[91]), .IN5(
          key[219]), .IN6(n6711), .QN(n3028));
   AOI222X1 U4783 (.IN1(n2484), .IN2(n7050), .IN3(n2481), .IN4(n7139), .IN5(n2483), .IN6(
          n7105), .QN(n3032));
   XNOR2X1 U4784 (.IN1(n3033), .IN2(n2960), .Q(n2483));
   XNOR2X1 U4785 (.IN1(n7593), .IN2(n3033), .Q(n2481));
   XNOR2X1 U4786 (.IN1(prev_key0_reg[90]), .IN2(n2220), .Q(n3033));
   XOR3X1 U4787 (.IN1(prev_key1_reg[90]), .IN2(prev_key1_reg[122]), .IN3(n7585), .Q(n2484)
          );
   AOI222X1 U4788 (.IN1(prev_key1_reg[90]), .IN2(n6950), .IN3(n7084), .IN4(key[90]), .IN5(
          key[218]), .IN6(n6709), .QN(n3031));
   AOI222X1 U4789 (.IN1(n2489), .IN2(n7050), .IN3(n2486), .IN4(n7139), .IN5(n2488), .IN6(
          n7105), .QN(n3035));
   XNOR2X1 U4790 (.IN1(n3036), .IN2(n2963), .Q(n2488));
   XNOR2X1 U4791 (.IN1(n7592), .IN2(n3036), .Q(n2486));
   XNOR2X1 U4792 (.IN1(prev_key0_reg[89]), .IN2(n2221), .Q(n3036));
   XOR3X1 U4793 (.IN1(prev_key1_reg[89]), .IN2(prev_key1_reg[121]), .IN3(n7584), .Q(n2489)
          );
   AOI222X1 U4794 (.IN1(prev_key1_reg[89]), .IN2(n6954), .IN3(n7084), .IN4(key[89]), .IN5(
          key[217]), .IN6(n6710), .QN(n3034));
   AOI222X1 U4795 (.IN1(n2494), .IN2(n7050), .IN3(n2491), .IN4(n7139), .IN5(n2493), .IN6(
          n7105), .QN(n3038));
   XNOR2X1 U4796 (.IN1(n3039), .IN2(n2966), .Q(n2493));
   XNOR2X1 U4797 (.IN1(n7591), .IN2(n3039), .Q(n2491));
   XNOR2X1 U4798 (.IN1(prev_key0_reg[88]), .IN2(n2222), .Q(n3039));
   XOR3X1 U4799 (.IN1(prev_key1_reg[88]), .IN2(prev_key1_reg[120]), .IN3(n7583), .Q(n2494)
          );
   AOI222X1 U4800 (.IN1(prev_key1_reg[88]), .IN2(n6951), .IN3(n7084), .IN4(key[88]), .IN5(
          key[216]), .IN6(n6709), .QN(n3037));
   AOI222X1 U4801 (.IN1(n2499), .IN2(n7051), .IN3(n2496), .IN4(n7139), .IN5(n2498), .IN6(
          n7105), .QN(n3041));
   XOR2X1 U4802 (.IN1(new_sboxw[15]), .IN2(n3042), .Q(n2498));
   XOR2X1 U4803 (.IN1(new_sboxw[23]), .IN2(n3042), .Q(n2496));
   XOR2X1 U4804 (.IN1(prev_key0_reg[87]), .IN2(prev_key0_reg[119]), .Q(n3042));
   XOR3X1 U4805 (.IN1(prev_key1_reg[87]), .IN2(prev_key1_reg[119]), .IN3(new_sboxw[15]), .
          Q(n2499));
   AOI222X1 U4806 (.IN1(prev_key1_reg[87]), .IN2(n6951), .IN3(n7084), .IN4(key[87]), .IN5(
          key[215]), .IN6(n6706), .QN(n3040));
   AOI222X1 U4807 (.IN1(n2504), .IN2(n7051), .IN3(n2501), .IN4(n7139), .IN5(n2503), .IN6(
          n7105), .QN(n3044));
   XOR2X1 U4808 (.IN1(new_sboxw[14]), .IN2(n3045), .Q(n2503));
   XOR2X1 U4810 (.IN1(prev_key0_reg[86]), .IN2(prev_key0_reg[118]), .Q(n3045));
   XOR3X1 U4811 (.IN1(prev_key1_reg[86]), .IN2(prev_key1_reg[118]), .IN3(new_sboxw[14]), .
          Q(n2504));
   AOI222X1 U4812 (.IN1(prev_key1_reg[86]), .IN2(n6952), .IN3(n7084), .IN4(key[86]), .IN5(
          key[214]), .IN6(n6705), .QN(n3043));
   AOI222X1 U4813 (.IN1(n2509), .IN2(n7051), .IN3(n2506), .IN4(n7139), .IN5(n2508), .IN6(
          n7105), .QN(n3047));
   XOR2X1 U4814 (.IN1(new_sboxw[13]), .IN2(n3048), .Q(n2508));
   XOR2X1 U4815 (.IN1(new_sboxw[21]), .IN2(n3048), .Q(n2506));
   XOR2X1 U4816 (.IN1(prev_key0_reg[85]), .IN2(prev_key0_reg[117]), .Q(n3048));
   XOR3X1 U4817 (.IN1(prev_key1_reg[85]), .IN2(prev_key1_reg[117]), .IN3(new_sboxw[13]), .
          Q(n2509));
   AOI222X1 U4818 (.IN1(prev_key1_reg[85]), .IN2(n6953), .IN3(n7084), .IN4(key[85]), .IN5(
          key[213]), .IN6(n6708), .QN(n3046));
   AOI222X1 U4819 (.IN1(n2514), .IN2(n7051), .IN3(n2511), .IN4(n7139), .IN5(n2513), .IN6(
          n7105), .QN(n3050));
   XOR2X1 U4820 (.IN1(new_sboxw[12]), .IN2(n3051), .Q(n2513));
   XOR2X1 U4821 (.IN1(new_sboxw[20]), .IN2(n3051), .Q(n2511));
   XOR2X1 U4822 (.IN1(prev_key0_reg[84]), .IN2(prev_key0_reg[116]), .Q(n3051));
   XOR3X1 U4823 (.IN1(prev_key1_reg[84]), .IN2(prev_key1_reg[116]), .IN3(new_sboxw[12]), .
          Q(n2514));
   AOI222X1 U4824 (.IN1(prev_key1_reg[84]), .IN2(n6954), .IN3(n7084), .IN4(key[84]), .IN5(
          key[212]), .IN6(n6707), .QN(n3049));
   AOI222X1 U4825 (.IN1(n2519), .IN2(n7051), .IN3(n2516), .IN4(n7140), .IN5(n2518), .IN6(
          n7104), .QN(n3053));
   XOR2X1 U4826 (.IN1(new_sboxw[11]), .IN2(n3054), .Q(n2518));
   XOR2X1 U4827 (.IN1(new_sboxw[19]), .IN2(n3054), .Q(n2516));
   XOR2X1 U4828 (.IN1(prev_key0_reg[83]), .IN2(prev_key0_reg[115]), .Q(n3054));
   XOR3X1 U4829 (.IN1(prev_key1_reg[83]), .IN2(prev_key1_reg[115]), .IN3(new_sboxw[11]), .
          Q(n2519));
   AOI222X1 U4830 (.IN1(prev_key1_reg[83]), .IN2(n6947), .IN3(n7084), .IN4(key[83]), .IN5(
          key[211]), .IN6(n6706), .QN(n3052));
   AOI222X1 U4831 (.IN1(n2524), .IN2(n7051), .IN3(n2521), .IN4(n7140), .IN5(n2523), .IN6(
          n7104), .QN(n3056));
   XOR2X1 U4832 (.IN1(new_sboxw[10]), .IN2(n3057), .Q(n2523));
   XOR2X1 U4833 (.IN1(new_sboxw[18]), .IN2(n3057), .Q(n2521));
   XOR2X1 U4834 (.IN1(prev_key0_reg[82]), .IN2(prev_key0_reg[114]), .Q(n3057));
   XOR3X1 U4835 (.IN1(prev_key1_reg[82]), .IN2(prev_key1_reg[114]), .IN3(new_sboxw[10]), .
          Q(n2524));
   AOI222X1 U4836 (.IN1(prev_key1_reg[82]), .IN2(n6946), .IN3(n7084), .IN4(key[82]), .IN5(
          key[210]), .IN6(n6705), .QN(n3055));
   AOI222X1 U4837 (.IN1(n2529), .IN2(n7051), .IN3(n2526), .IN4(n7140), .IN5(n2528), .IN6(
          n7104), .QN(n3059));
   XOR2X1 U4838 (.IN1(new_sboxw[9]), .IN2(n3060), .Q(n2528));
   XOR2X1 U4839 (.IN1(new_sboxw[17]), .IN2(n3060), .Q(n2526));
   XOR2X1 U4840 (.IN1(prev_key0_reg[81]), .IN2(prev_key0_reg[113]), .Q(n3060));
   XOR3X1 U4841 (.IN1(prev_key1_reg[81]), .IN2(prev_key1_reg[113]), .IN3(new_sboxw[9]), .Q(
          n2529));
   AOI222X1 U4842 (.IN1(prev_key1_reg[81]), .IN2(n6955), .IN3(n7084), .IN4(key[81]), .IN5(
          key[209]), .IN6(n6704), .QN(n3058));
   AOI222X1 U4843 (.IN1(n2534), .IN2(n7051), .IN3(n2531), .IN4(n7140), .IN5(n2533), .IN6(
          n7104), .QN(n3062));
   XOR2X1 U4844 (.IN1(new_sboxw[8]), .IN2(n3063), .Q(n2533));
   XOR2X1 U4845 (.IN1(new_sboxw[16]), .IN2(n3063), .Q(n2531));
   XOR2X1 U4846 (.IN1(prev_key0_reg[80]), .IN2(prev_key0_reg[112]), .Q(n3063));
   XOR3X1 U4847 (.IN1(prev_key1_reg[80]), .IN2(prev_key1_reg[112]), .IN3(new_sboxw[8]), .Q(
          n2534));
   AOI222X1 U4848 (.IN1(prev_key1_reg[80]), .IN2(n6947), .IN3(n7085), .IN4(key[80]), .IN5(
          key[208]), .IN6(n6703), .QN(n3061));
   AOI222X1 U4849 (.IN1(n2539), .IN2(n7051), .IN3(n2536), .IN4(n7140), .IN5(n2538), .IN6(
          n7104), .QN(n3065));
   XOR2X1 U4851 (.IN1(new_sboxw[15]), .IN2(n3066), .Q(n2536));
   XOR2X1 U4852 (.IN1(prev_key0_reg[79]), .IN2(prev_key0_reg[111]), .Q(n3066));
   AOI222X1 U4854 (.IN1(prev_key1_reg[79]), .IN2(n6953), .IN3(n7085), .IN4(key[79]), .IN5(
          key[207]), .IN6(n6711), .QN(n3064));
   AOI222X1 U4855 (.IN1(n2544), .IN2(n7051), .IN3(n2541), .IN4(n7140), .IN5(n2543), .IN6(
          n7104), .QN(n3068));
   XOR2X1 U4856 (.IN1(new_sboxw[6]), .IN2(n3069), .Q(n2543));
   XOR2X1 U4857 (.IN1(new_sboxw[14]), .IN2(n3069), .Q(n2541));
   XOR2X1 U4858 (.IN1(prev_key0_reg[78]), .IN2(prev_key0_reg[110]), .Q(n3069));
   XOR3X1 U4859 (.IN1(prev_key1_reg[78]), .IN2(prev_key1_reg[110]), .IN3(new_sboxw[6]), .Q(
          n2544));
   AOI222X1 U4860 (.IN1(prev_key1_reg[78]), .IN2(n6954), .IN3(n7085), .IN4(key[78]), .IN5(
          key[206]), .IN6(n6708), .QN(n3067));
   AOI222X1 U4861 (.IN1(n2549), .IN2(n7051), .IN3(n2546), .IN4(n7140), .IN5(n2548), .IN6(
          n7104), .QN(n3071));
   XOR2X1 U4863 (.IN1(new_sboxw[13]), .IN2(n3072), .Q(n2546));
   XOR2X1 U4864 (.IN1(prev_key0_reg[77]), .IN2(prev_key0_reg[109]), .Q(n3072));
   AOI222X1 U4866 (.IN1(prev_key1_reg[77]), .IN2(n6944), .IN3(n7085), .IN4(key[77]), .IN5(
          key[205]), .IN6(n6704), .QN(n3070));
   AOI222X1 U4867 (.IN1(n2554), .IN2(n7051), .IN3(n2551), .IN4(n7140), .IN5(n2553), .IN6(
          n7104), .QN(n3074));
   XOR2X1 U4868 (.IN1(new_sboxw[4]), .IN2(n3075), .Q(n2553));
   XOR2X1 U4869 (.IN1(new_sboxw[12]), .IN2(n3075), .Q(n2551));
   XOR2X1 U4870 (.IN1(prev_key0_reg[76]), .IN2(prev_key0_reg[108]), .Q(n3075));
   XOR3X1 U4871 (.IN1(prev_key1_reg[76]), .IN2(prev_key1_reg[108]), .IN3(new_sboxw[4]), .Q(
          n2554));
   AOI222X1 U4872 (.IN1(prev_key1_reg[76]), .IN2(n6947), .IN3(n7085), .IN4(key[76]), .IN5(
          key[204]), .IN6(n6703), .QN(n3073));
   AOI222X1 U4873 (.IN1(n2559), .IN2(n7051), .IN3(n2556), .IN4(n7140), .IN5(n2558), .IN6(
          n7104), .QN(n3077));
   XOR2X1 U4874 (.IN1(new_sboxw[3]), .IN2(n3078), .Q(n2558));
   XOR2X1 U4875 (.IN1(new_sboxw[11]), .IN2(n3078), .Q(n2556));
   XOR2X1 U4876 (.IN1(prev_key0_reg[75]), .IN2(prev_key0_reg[107]), .Q(n3078));
   XOR3X1 U4877 (.IN1(prev_key1_reg[75]), .IN2(prev_key1_reg[107]), .IN3(new_sboxw[3]), .Q(
          n2559));
   AOI222X1 U4878 (.IN1(prev_key1_reg[75]), .IN2(n6951), .IN3(n7085), .IN4(key[75]), .IN5(
          key[203]), .IN6(n6710), .QN(n3076));
   AOI222X1 U4879 (.IN1(n2564), .IN2(n7051), .IN3(n2561), .IN4(n7140), .IN5(n2563), .IN6(
          n7104), .QN(n3080));
   XOR2X1 U4881 (.IN1(new_sboxw[10]), .IN2(n3081), .Q(n2561));
   XOR2X1 U4882 (.IN1(prev_key0_reg[74]), .IN2(prev_key0_reg[106]), .Q(n3081));
   AOI222X1 U4884 (.IN1(prev_key1_reg[74]), .IN2(n6952), .IN3(n7085), .IN4(key[74]), .IN5(
          key[202]), .IN6(n6709), .QN(n3079));
   AOI222X1 U4885 (.IN1(n2569), .IN2(n7051), .IN3(n2566), .IN4(n7140), .IN5(n2568), .IN6(
          n7104), .QN(n3083));
   XOR2X1 U4887 (.IN1(new_sboxw[9]), .IN2(n3084), .Q(n2566));
   XOR2X1 U4888 (.IN1(prev_key0_reg[73]), .IN2(prev_key0_reg[105]), .Q(n3084));
   AOI222X1 U4890 (.IN1(prev_key1_reg[73]), .IN2(n6952), .IN3(n7085), .IN4(key[73]), .IN5(
          key[201]), .IN6(n6708), .QN(n3082));
   AOI222X1 U4891 (.IN1(n2574), .IN2(n7051), .IN3(n2571), .IN4(n7140), .IN5(n2573), .IN6(
          n7104), .QN(n3086));
   XOR2X1 U4892 (.IN1(new_sboxw[0]), .IN2(n3087), .Q(n2573));
   XOR2X1 U4893 (.IN1(new_sboxw[8]), .IN2(n3087), .Q(n2571));
   XOR2X1 U4894 (.IN1(prev_key0_reg[72]), .IN2(prev_key0_reg[104]), .Q(n3087));
   XOR3X1 U4895 (.IN1(prev_key1_reg[72]), .IN2(prev_key1_reg[104]), .IN3(new_sboxw[0]), .Q(
          n2574));
   AOI222X1 U4896 (.IN1(prev_key1_reg[72]), .IN2(n6953), .IN3(n7085), .IN4(key[72]), .IN5(
          key[200]), .IN6(n6707), .QN(n3085));
   AOI222X1 U4897 (.IN1(n2579), .IN2(n7051), .IN3(n2576), .IN4(n7140), .IN5(n2578), .IN6(
          n7103), .QN(n3089));
   XOR2X1 U4898 (.IN1(new_sboxw[31]), .IN2(n3090), .Q(n2578));
   XOR2X1 U4900 (.IN1(prev_key0_reg[71]), .IN2(prev_key0_reg[103]), .Q(n3090));
   XOR3X1 U4901 (.IN1(prev_key1_reg[71]), .IN2(prev_key1_reg[103]), .IN3(new_sboxw[31]), .
          Q(n2579));
   AOI222X1 U4902 (.IN1(prev_key1_reg[71]), .IN2(n6954), .IN3(n7085), .IN4(key[71]), .IN5(
          key[199]), .IN6(n6706), .QN(n3088));
   AOI222X1 U4903 (.IN1(n2584), .IN2(n7052), .IN3(n2581), .IN4(n7141), .IN5(n2583), .IN6(
          n7103), .QN(n3092));
   XOR2X1 U4904 (.IN1(new_sboxw[30]), .IN2(n3093), .Q(n2583));
   XOR2X1 U4905 (.IN1(new_sboxw[6]), .IN2(n3093), .Q(n2581));
   XOR2X1 U4906 (.IN1(prev_key0_reg[70]), .IN2(prev_key0_reg[102]), .Q(n3093));
   XOR3X1 U4907 (.IN1(prev_key1_reg[70]), .IN2(prev_key1_reg[102]), .IN3(new_sboxw[30]), .
          Q(n2584));
   AOI222X1 U4908 (.IN1(prev_key1_reg[70]), .IN2(n6945), .IN3(n7085), .IN4(key[70]), .IN5(
          key[198]), .IN6(n6705), .QN(n3091));
   AOI222X1 U4909 (.IN1(n2589), .IN2(n7052), .IN3(n2586), .IN4(n7141), .IN5(n2588), .IN6(
          n7103), .QN(n3095));
   XOR2X1 U4910 (.IN1(new_sboxw[29]), .IN2(n3096), .Q(n2588));
   XOR2X1 U4912 (.IN1(prev_key0_reg[69]), .IN2(prev_key0_reg[101]), .Q(n3096));
   XOR3X1 U4913 (.IN1(prev_key1_reg[69]), .IN2(prev_key1_reg[101]), .IN3(new_sboxw[29]), .
          Q(n2589));
   AOI222X1 U4914 (.IN1(prev_key1_reg[69]), .IN2(n6946), .IN3(n7085), .IN4(key[69]), .IN5(
          key[197]), .IN6(n6704), .QN(n3094));
   AOI222X1 U4915 (.IN1(n2594), .IN2(n7052), .IN3(n2591), .IN4(n7141), .IN5(n2593), .IN6(
          n7103), .QN(n3098));
   XOR2X1 U4916 (.IN1(new_sboxw[28]), .IN2(n3099), .Q(n2593));
   XOR2X1 U4917 (.IN1(new_sboxw[4]), .IN2(n3099), .Q(n2591));
   XOR2X1 U4918 (.IN1(prev_key0_reg[68]), .IN2(prev_key0_reg[100]), .Q(n3099));
   XOR3X1 U4919 (.IN1(prev_key1_reg[68]), .IN2(prev_key1_reg[100]), .IN3(new_sboxw[28]), .
          Q(n2594));
   AOI222X1 U4920 (.IN1(prev_key1_reg[68]), .IN2(n6947), .IN3(n7085), .IN4(key[68]), .IN5(
          key[196]), .IN6(n6703), .QN(n3097));
   AOI222X1 U4921 (.IN1(n2599), .IN2(n7052), .IN3(n2596), .IN4(n7141), .IN5(n2598), .IN6(
          n7103), .QN(n3101));
   XOR2X1 U4922 (.IN1(new_sboxw[27]), .IN2(n3102), .Q(n2598));
   XOR2X1 U4923 (.IN1(new_sboxw[3]), .IN2(n3102), .Q(n2596));
   XOR2X1 U4924 (.IN1(prev_key0_reg[67]), .IN2(prev_key0_reg[99]), .Q(n3102));
   XOR3X1 U4925 (.IN1(prev_key1_reg[99]), .IN2(prev_key1_reg[67]), .IN3(new_sboxw[27]), .Q(
          n2599));
   AOI222X1 U4926 (.IN1(prev_key1_reg[67]), .IN2(n6948), .IN3(n7085), .IN4(key[67]), .IN5(
          key[195]), .IN6(n6711), .QN(n3100));
   AOI222X1 U4927 (.IN1(n2604), .IN2(n7052), .IN3(n2601), .IN4(n7141), .IN5(n2603), .IN6(
          n7103), .QN(n3104));
   XOR2X1 U4928 (.IN1(new_sboxw[26]), .IN2(n3105), .Q(n2603));
   XOR2X1 U4930 (.IN1(prev_key0_reg[66]), .IN2(prev_key0_reg[98]), .Q(n3105));
   XOR3X1 U4931 (.IN1(prev_key1_reg[98]), .IN2(prev_key1_reg[66]), .IN3(new_sboxw[26]), .Q(
          n2604));
   AOI222X1 U4932 (.IN1(prev_key1_reg[66]), .IN2(n6949), .IN3(n7086), .IN4(key[66]), .IN5(
          key[194]), .IN6(n6711), .QN(n3103));
   AOI222X1 U4933 (.IN1(n2609), .IN2(n7052), .IN3(n2606), .IN4(n7141), .IN5(n2608), .IN6(
          n7103), .QN(n3107));
   XOR2X1 U4934 (.IN1(new_sboxw[25]), .IN2(n3108), .Q(n2608));
   XOR2X1 U4936 (.IN1(prev_key0_reg[65]), .IN2(prev_key0_reg[97]), .Q(n3108));
   XOR3X1 U4937 (.IN1(prev_key1_reg[97]), .IN2(prev_key1_reg[65]), .IN3(new_sboxw[25]), .Q(
          n2609));
   AOI222X1 U4938 (.IN1(prev_key1_reg[65]), .IN2(n6954), .IN3(n7086), .IN4(key[65]), .IN5(
          key[193]), .IN6(n6711), .QN(n3106));
   AOI222X1 U4939 (.IN1(n2614), .IN2(n7052), .IN3(n2611), .IN4(n7141), .IN5(n2613), .IN6(
          n7103), .QN(n3110));
   XOR2X1 U4940 (.IN1(new_sboxw[24]), .IN2(n3111), .Q(n2613));
   XOR2X1 U4941 (.IN1(new_sboxw[0]), .IN2(n3111), .Q(n2611));
   XOR2X1 U4942 (.IN1(prev_key0_reg[64]), .IN2(prev_key0_reg[96]), .Q(n3111));
   XOR3X1 U4943 (.IN1(prev_key1_reg[96]), .IN2(prev_key1_reg[64]), .IN3(new_sboxw[24]), .Q(
          n2614));
   AOI222X1 U4944 (.IN1(prev_key1_reg[64]), .IN2(n6950), .IN3(n7086), .IN4(key[64]), .IN5(
          key[192]), .IN6(n6711), .QN(n3109));
   AOI222X1 U4945 (.IN1(n2619), .IN2(n7052), .IN3(n2616), .IN4(n7141), .IN5(n2618), .IN6(
          n7103), .QN(n3113));
   XOR2X1 U4946 (.IN1(n3114), .IN2(n7590), .Q(n2618));
   XOR2X1 U4947 (.IN1(n3114), .IN2(n7598), .Q(n2616));
   XNOR3X1 U4948 (.IN1(prev_key0_reg[95]), .IN2(prev_key0_reg[63]), .IN3(
          prev_key0_reg[127]), .Q(n3114));
   XNOR3X1 U4949 (.IN1(prev_key1_reg[95]), .IN2(prev_key1_reg[63]), .IN3(n3115), .Q(n2619)
          );
   XNOR2X1 U4950 (.IN1(prev_key1_reg[127]), .IN2(n3018), .Q(n3115));
   AOI222X1 U4951 (.IN1(prev_key1_reg[63]), .IN2(n6951), .IN3(n7086), .IN4(key[63]), .IN5(
          key[191]), .IN6(n6710), .QN(n3112));
   AOI222X1 U4952 (.IN1(n2624), .IN2(n7052), .IN3(n2621), .IN4(n7141), .IN5(n2623), .IN6(
          n7103), .QN(n3117));
   XOR2X1 U4953 (.IN1(n3118), .IN2(n2948), .Q(n2623));
   XOR2X1 U4954 (.IN1(n3118), .IN2(n7597), .Q(n2621));
   XNOR3X1 U4955 (.IN1(prev_key0_reg[94]), .IN2(prev_key0_reg[62]), .IN3(
          prev_key0_reg[126]), .Q(n3118));
   XNOR3X1 U4956 (.IN1(prev_key1_reg[94]), .IN2(prev_key1_reg[62]), .IN3(n3119), .Q(n2624)
          );
   XNOR2X1 U4957 (.IN1(prev_key1_reg[126]), .IN2(n7589), .Q(n3119));
   AOI222X1 U4958 (.IN1(prev_key1_reg[62]), .IN2(n6952), .IN3(n7086), .IN4(key[62]), .IN5(
          key[190]), .IN6(n6709), .QN(n3116));
   AOI222X1 U4959 (.IN1(n2629), .IN2(n7052), .IN3(n2626), .IN4(n7141), .IN5(n2628), .IN6(
          n7103), .QN(n3121));
   XOR2X1 U4960 (.IN1(n3122), .IN2(n2951), .Q(n2628));
   XOR2X1 U4961 (.IN1(n3122), .IN2(n7596), .Q(n2626));
   XNOR3X1 U4962 (.IN1(prev_key0_reg[93]), .IN2(prev_key0_reg[61]), .IN3(
          prev_key0_reg[125]), .Q(n3122));
   XNOR3X1 U4963 (.IN1(prev_key1_reg[93]), .IN2(prev_key1_reg[61]), .IN3(n3123), .Q(n2629)
          );
   XNOR2X1 U4964 (.IN1(prev_key1_reg[125]), .IN2(n7588), .Q(n3123));
   AOI222X1 U4965 (.IN1(prev_key1_reg[61]), .IN2(n6953), .IN3(n7086), .IN4(key[61]), .IN5(
          key[189]), .IN6(n6708), .QN(n3120));
   AOI222X1 U4966 (.IN1(n2634), .IN2(n7052), .IN3(n2631), .IN4(n7141), .IN5(n2633), .IN6(
          n7103), .QN(n3125));
   XOR2X1 U4967 (.IN1(n3126), .IN2(n2954), .Q(n2633));
   XOR2X1 U4968 (.IN1(n3126), .IN2(n7595), .Q(n2631));
   XNOR3X1 U4969 (.IN1(prev_key0_reg[92]), .IN2(prev_key0_reg[60]), .IN3(
          prev_key0_reg[124]), .Q(n3126));
   XNOR3X1 U4970 (.IN1(prev_key1_reg[92]), .IN2(prev_key1_reg[60]), .IN3(n3127), .Q(n2634)
          );
   XNOR2X1 U4971 (.IN1(prev_key1_reg[124]), .IN2(n7587), .Q(n3127));
   AOI222X1 U4972 (.IN1(prev_key1_reg[60]), .IN2(n6954), .IN3(n7086), .IN4(key[60]), .IN5(
          key[188]), .IN6(n6707), .QN(n3124));
   AOI222X1 U4973 (.IN1(n2639), .IN2(n7052), .IN3(n2636), .IN4(n7141), .IN5(n2638), .IN6(
          n7102), .QN(n3129));
   XOR2X1 U4974 (.IN1(n3130), .IN2(n2957), .Q(n2638));
   XOR2X1 U4975 (.IN1(n3130), .IN2(n7594), .Q(n2636));
   XNOR3X1 U4976 (.IN1(prev_key0_reg[91]), .IN2(prev_key0_reg[59]), .IN3(
          prev_key0_reg[123]), .Q(n3130));
   XNOR3X1 U4977 (.IN1(prev_key1_reg[91]), .IN2(prev_key1_reg[59]), .IN3(n3131), .Q(n2639)
          );
   XNOR2X1 U4978 (.IN1(prev_key1_reg[123]), .IN2(n7586), .Q(n3131));
   AOI222X1 U4979 (.IN1(prev_key1_reg[59]), .IN2(n6948), .IN3(n7086), .IN4(key[59]), .IN5(
          key[187]), .IN6(n6706), .QN(n3128));
   AOI222X1 U4980 (.IN1(n2644), .IN2(n7052), .IN3(n2641), .IN4(n7141), .IN5(n2643), .IN6(
          n7102), .QN(n3133));
   XOR2X1 U4981 (.IN1(n3134), .IN2(n2960), .Q(n2643));
   XOR2X1 U4982 (.IN1(n3134), .IN2(n7593), .Q(n2641));
   XNOR3X1 U4983 (.IN1(prev_key0_reg[90]), .IN2(prev_key0_reg[58]), .IN3(
          prev_key0_reg[122]), .Q(n3134));
   XNOR3X1 U4984 (.IN1(prev_key1_reg[90]), .IN2(prev_key1_reg[58]), .IN3(n3135), .Q(n2644)
          );
   XNOR2X1 U4985 (.IN1(prev_key1_reg[122]), .IN2(n7585), .Q(n3135));
   AOI222X1 U4986 (.IN1(prev_key1_reg[58]), .IN2(n6948), .IN3(n7086), .IN4(key[58]), .IN5(
          key[186]), .IN6(n6705), .QN(n3132));
   AOI222X1 U4987 (.IN1(n2649), .IN2(n7052), .IN3(n2646), .IN4(n7142), .IN5(n2648), .IN6(
          n7102), .QN(n3137));
   XOR2X1 U4988 (.IN1(n3138), .IN2(n2963), .Q(n2648));
   XOR2X1 U4989 (.IN1(n3138), .IN2(n7592), .Q(n2646));
   XNOR3X1 U4990 (.IN1(prev_key0_reg[89]), .IN2(prev_key0_reg[57]), .IN3(
          prev_key0_reg[121]), .Q(n3138));
   XNOR3X1 U4991 (.IN1(prev_key1_reg[89]), .IN2(prev_key1_reg[57]), .IN3(n3139), .Q(n2649)
          );
   XNOR2X1 U4992 (.IN1(prev_key1_reg[121]), .IN2(n7584), .Q(n3139));
   AOI222X1 U4993 (.IN1(prev_key1_reg[57]), .IN2(n6953), .IN3(n7086), .IN4(key[57]), .IN5(
          key[185]), .IN6(n6710), .QN(n3136));
   AOI222X1 U4994 (.IN1(n2654), .IN2(n7052), .IN3(n2651), .IN4(n7142), .IN5(n2653), .IN6(
          n7102), .QN(n3141));
   XOR2X1 U4995 (.IN1(n3142), .IN2(n2966), .Q(n2653));
   XOR2X1 U4996 (.IN1(n3142), .IN2(n7591), .Q(n2651));
   XNOR3X1 U4997 (.IN1(prev_key0_reg[88]), .IN2(prev_key0_reg[56]), .IN3(
          prev_key0_reg[120]), .Q(n3142));
   AOI222X1 U5000 (.IN1(prev_key1_reg[56]), .IN2(n6954), .IN3(n7086), .IN4(key[56]), .IN5(
          key[184]), .IN6(n6709), .QN(n3140));
   AOI222X1 U5001 (.IN1(n2659), .IN2(n7052), .IN3(n2656), .IN4(n7142), .IN5(n2658), .IN6(
          n7102), .QN(n3145));
   XOR2X1 U5002 (.IN1(n3146), .IN2(n7611), .Q(n2658));
   XNOR2X1 U5003 (.IN1(n3146), .IN2(new_sboxw[23]), .Q(n2656));
   XNOR3X1 U5004 (.IN1(prev_key0_reg[87]), .IN2(prev_key0_reg[55]), .IN3(
          prev_key0_reg[119]), .Q(n3146));
   XNOR3X1 U5005 (.IN1(prev_key1_reg[119]), .IN2(new_sboxw[15]), .IN3(n3147), .Q(n2659));
   XNOR2X1 U5006 (.IN1(prev_key1_reg[55]), .IN2(prev_key1_reg[87]), .Q(n3147));
   AOI222X1 U5007 (.IN1(prev_key1_reg[55]), .IN2(n6949), .IN3(n7086), .IN4(key[55]), .IN5(
          key[183]), .IN6(n6704), .QN(n3144));
   AOI222X1 U5008 (.IN1(n2664), .IN2(n7052), .IN3(n2661), .IN4(n7142), .IN5(n2663), .IN6(
          n7102), .QN(n3149));
   XOR2X1 U5009 (.IN1(n3150), .IN2(n6700), .Q(n2663));
   XOR2X1 U5010 (.IN1(n3150), .IN2(n7605), .Q(n2661));
   XNOR3X1 U5011 (.IN1(prev_key0_reg[86]), .IN2(prev_key0_reg[54]), .IN3(
          prev_key0_reg[118]), .Q(n3150));
   XNOR3X1 U5012 (.IN1(prev_key1_reg[118]), .IN2(new_sboxw[14]), .IN3(n3151), .Q(n2664));
   XNOR2X1 U5013 (.IN1(prev_key1_reg[54]), .IN2(prev_key1_reg[86]), .Q(n3151));
   AOI222X1 U5014 (.IN1(prev_key1_reg[54]), .IN2(n6948), .IN3(n7086), .IN4(key[54]), .IN5(
          key[182]), .IN6(n6703), .QN(n3148));
   AOI222X1 U5015 (.IN1(n2669), .IN2(n7053), .IN3(n2666), .IN4(n7142), .IN5(n2668), .IN6(
          n7102), .QN(n3153));
   XOR2X1 U5016 (.IN1(n3154), .IN2(n7609), .Q(n2668));
   XOR2X1 U5017 (.IN1(n3154), .IN2(n7604), .Q(n2666));
   XNOR3X1 U5018 (.IN1(prev_key0_reg[85]), .IN2(prev_key0_reg[53]), .IN3(
          prev_key0_reg[117]), .Q(n3154));
   XNOR3X1 U5019 (.IN1(prev_key1_reg[117]), .IN2(new_sboxw[13]), .IN3(n3155), .Q(n2669));
   XNOR2X1 U5020 (.IN1(prev_key1_reg[53]), .IN2(prev_key1_reg[85]), .Q(n3155));
   AOI222X1 U5021 (.IN1(prev_key1_reg[53]), .IN2(n6955), .IN3(n7086), .IN4(key[53]), .IN5(
          key[181]), .IN6(n6711), .QN(n3152));
   AOI222X1 U5022 (.IN1(n2674), .IN2(n7053), .IN3(n2671), .IN4(n7142), .IN5(n2673), .IN6(
          n7102), .QN(n3157));
   XOR2X1 U5023 (.IN1(n3158), .IN2(n7608), .Q(n2673));
   XOR2X1 U5024 (.IN1(n3158), .IN2(n7603), .Q(n2671));
   XNOR3X1 U5025 (.IN1(prev_key0_reg[84]), .IN2(prev_key0_reg[52]), .IN3(
          prev_key0_reg[116]), .Q(n3158));
   XNOR3X1 U5026 (.IN1(prev_key1_reg[116]), .IN2(new_sboxw[12]), .IN3(n3159), .Q(n2674));
   XNOR2X1 U5027 (.IN1(prev_key1_reg[52]), .IN2(prev_key1_reg[84]), .Q(n3159));
   AOI222X1 U5028 (.IN1(prev_key1_reg[52]), .IN2(n6949), .IN3(n7087), .IN4(key[52]), .IN5(
          key[180]), .IN6(n2945), .QN(n3156));
   AOI222X1 U5029 (.IN1(n2679), .IN2(n7053), .IN3(n2676), .IN4(n7142), .IN5(n2678), .IN6(
          n7102), .QN(n3161));
   XOR2X1 U5030 (.IN1(n3162), .IN2(n7607), .Q(n2678));
   XOR2X1 U5031 (.IN1(n3162), .IN2(n7602), .Q(n2676));
   XNOR3X1 U5032 (.IN1(prev_key0_reg[83]), .IN2(prev_key0_reg[51]), .IN3(
          prev_key0_reg[115]), .Q(n3162));
   XNOR3X1 U5033 (.IN1(prev_key1_reg[115]), .IN2(new_sboxw[11]), .IN3(n3163), .Q(n2679));
   XNOR2X1 U5034 (.IN1(prev_key1_reg[51]), .IN2(prev_key1_reg[83]), .Q(n3163));
   AOI222X1 U5035 (.IN1(prev_key1_reg[51]), .IN2(n6955), .IN3(n7087), .IN4(key[51]), .IN5(
          key[179]), .IN6(n6710), .QN(n3160));
   AOI222X1 U5036 (.IN1(n2684), .IN2(n7053), .IN3(n2681), .IN4(n7142), .IN5(n2683), .IN6(
          n7102), .QN(n3165));
   XOR2X1 U5037 (.IN1(n3166), .IN2(n7606), .Q(n2683));
   XOR2X1 U5038 (.IN1(n3166), .IN2(n7601), .Q(n2681));
   XNOR3X1 U5039 (.IN1(prev_key0_reg[82]), .IN2(prev_key0_reg[50]), .IN3(
          prev_key0_reg[114]), .Q(n3166));
   XNOR3X1 U5040 (.IN1(prev_key1_reg[114]), .IN2(new_sboxw[10]), .IN3(n3167), .Q(n2684));
   XNOR2X1 U5041 (.IN1(prev_key1_reg[50]), .IN2(prev_key1_reg[82]), .Q(n3167));
   AOI222X1 U5042 (.IN1(prev_key1_reg[50]), .IN2(n6955), .IN3(n7087), .IN4(key[50]), .IN5(
          key[178]), .IN6(n6709), .QN(n3164));
   AOI222X1 U5043 (.IN1(n2689), .IN2(n7053), .IN3(n2686), .IN4(n7142), .IN5(n2688), .IN6(
          n7102), .QN(n3169));
   XOR2X1 U5044 (.IN1(n3170), .IN2(n7613), .Q(n2688));
   XOR2X1 U5045 (.IN1(n3170), .IN2(n7600), .Q(n2686));
   XNOR3X1 U5046 (.IN1(prev_key0_reg[81]), .IN2(prev_key0_reg[49]), .IN3(
          prev_key0_reg[113]), .Q(n3170));
   XNOR3X1 U5047 (.IN1(prev_key1_reg[113]), .IN2(new_sboxw[9]), .IN3(n3171), .Q(n2689));
   XNOR2X1 U5048 (.IN1(prev_key1_reg[49]), .IN2(prev_key1_reg[81]), .Q(n3171));
   AOI222X1 U5049 (.IN1(prev_key1_reg[49]), .IN2(n6953), .IN3(n7087), .IN4(key[49]), .IN5(
          key[177]), .IN6(n6708), .QN(n3168));
   AOI222X1 U5050 (.IN1(n2694), .IN2(n7053), .IN3(n2691), .IN4(n7142), .IN5(n2693), .IN6(
          n7102), .QN(n3173));
   XOR2X1 U5051 (.IN1(n3174), .IN2(n7612), .Q(n2693));
   XOR2X1 U5052 (.IN1(n3174), .IN2(n7599), .Q(n2691));
   XNOR3X1 U5053 (.IN1(prev_key0_reg[80]), .IN2(prev_key0_reg[48]), .IN3(
          prev_key0_reg[112]), .Q(n3174));
   XNOR3X1 U5054 (.IN1(prev_key1_reg[112]), .IN2(new_sboxw[8]), .IN3(n3175), .Q(n2694));
   XNOR2X1 U5055 (.IN1(prev_key1_reg[48]), .IN2(prev_key1_reg[80]), .Q(n3175));
   AOI222X1 U5056 (.IN1(prev_key1_reg[48]), .IN2(n6947), .IN3(n7087), .IN4(key[48]), .IN5(
          key[176]), .IN6(n6707), .QN(n3172));
   AOI222X1 U5057 (.IN1(n2699), .IN2(n7053), .IN3(n2696), .IN4(n7142), .IN5(n2698), .IN6(
          n7101), .QN(n3177));
   XOR2X1 U5058 (.IN1(n3178), .IN2(n7621), .Q(n2698));
   XOR2X1 U5059 (.IN1(n3178), .IN2(n7611), .Q(n2696));
   XNOR3X1 U5060 (.IN1(prev_key0_reg[79]), .IN2(prev_key0_reg[47]), .IN3(
          prev_key0_reg[111]), .Q(n3178));
   XNOR3X1 U5061 (.IN1(prev_key1_reg[111]), .IN2(new_sboxw[7]), .IN3(n3179), .Q(n2699));
   XNOR2X1 U5062 (.IN1(prev_key1_reg[47]), .IN2(prev_key1_reg[79]), .Q(n3179));
   AOI222X1 U5063 (.IN1(prev_key1_reg[47]), .IN2(n6944), .IN3(n7087), .IN4(key[47]), .IN5(
          key[175]), .IN6(n6708), .QN(n3176));
   AOI222X1 U5064 (.IN1(n2704), .IN2(n7053), .IN3(n2701), .IN4(n7142), .IN5(n2703), .IN6(
          n7101), .QN(n3181));
   XOR2X1 U5065 (.IN1(n3182), .IN2(n7620), .Q(n2703));
   XOR2X1 U5066 (.IN1(n3182), .IN2(n6700), .Q(n2701));
   XNOR3X1 U5067 (.IN1(prev_key0_reg[78]), .IN2(prev_key0_reg[46]), .IN3(
          prev_key0_reg[110]), .Q(n3182));
   XNOR3X1 U5068 (.IN1(prev_key1_reg[110]), .IN2(new_sboxw[6]), .IN3(n3183), .Q(n2704));
   XNOR2X1 U5069 (.IN1(prev_key1_reg[46]), .IN2(prev_key1_reg[78]), .Q(n3183));
   AOI222X1 U5070 (.IN1(prev_key1_reg[46]), .IN2(n6945), .IN3(n7087), .IN4(key[46]), .IN5(
          key[174]), .IN6(n6707), .QN(n3180));
   AOI222X1 U5071 (.IN1(n2709), .IN2(n7053), .IN3(n2706), .IN4(n7142), .IN5(n2708), .IN6(
          n7101), .QN(n3185));
   XOR2X1 U5072 (.IN1(n3186), .IN2(n7619), .Q(n2708));
   XOR2X1 U5073 (.IN1(n3186), .IN2(n7609), .Q(n2706));
   XNOR3X1 U5074 (.IN1(prev_key0_reg[77]), .IN2(prev_key0_reg[45]), .IN3(
          prev_key0_reg[109]), .Q(n3186));
   AOI222X1 U5077 (.IN1(prev_key1_reg[45]), .IN2(n6946), .IN3(n7087), .IN4(key[45]), .IN5(
          key[173]), .IN6(n6706), .QN(n3184));
   AOI222X1 U5078 (.IN1(n2714), .IN2(n7053), .IN3(n2711), .IN4(n7143), .IN5(n2713), .IN6(
          n7101), .QN(n3189));
   XOR2X1 U5079 (.IN1(n3190), .IN2(n7618), .Q(n2713));
   XOR2X1 U5080 (.IN1(n3190), .IN2(n7608), .Q(n2711));
   XNOR3X1 U5081 (.IN1(prev_key0_reg[76]), .IN2(prev_key0_reg[44]), .IN3(
          prev_key0_reg[108]), .Q(n3190));
   XNOR3X1 U5082 (.IN1(prev_key1_reg[108]), .IN2(new_sboxw[4]), .IN3(n3191), .Q(n2714));
   XNOR2X1 U5083 (.IN1(prev_key1_reg[44]), .IN2(prev_key1_reg[76]), .Q(n3191));
   AOI222X1 U5084 (.IN1(prev_key1_reg[44]), .IN2(n6947), .IN3(n7087), .IN4(key[44]), .IN5(
          key[172]), .IN6(n6705), .QN(n3188));
   AOI222X1 U5085 (.IN1(n2719), .IN2(n7053), .IN3(n2716), .IN4(n7143), .IN5(n2718), .IN6(
          n7101), .QN(n3193));
   XOR2X1 U5086 (.IN1(n3194), .IN2(n7617), .Q(n2718));
   XOR2X1 U5087 (.IN1(n3194), .IN2(n7607), .Q(n2716));
   XNOR3X1 U5088 (.IN1(prev_key0_reg[75]), .IN2(prev_key0_reg[43]), .IN3(
          prev_key0_reg[107]), .Q(n3194));
   XNOR3X1 U5089 (.IN1(prev_key1_reg[107]), .IN2(new_sboxw[3]), .IN3(n3195), .Q(n2719));
   XNOR2X1 U5090 (.IN1(prev_key1_reg[43]), .IN2(prev_key1_reg[75]), .Q(n3195));
   AOI222X1 U5091 (.IN1(prev_key1_reg[43]), .IN2(n6948), .IN3(n7087), .IN4(key[43]), .IN5(
          key[171]), .IN6(n6704), .QN(n3192));
   AOI222X1 U5092 (.IN1(n2724), .IN2(n7053), .IN3(n2721), .IN4(n7143), .IN5(n2723), .IN6(
          n7101), .QN(n3197));
   XOR2X1 U5093 (.IN1(n3198), .IN2(n7616), .Q(n2723));
   XOR2X1 U5094 (.IN1(n3198), .IN2(n7606), .Q(n2721));
   XNOR3X1 U5095 (.IN1(prev_key0_reg[74]), .IN2(prev_key0_reg[42]), .IN3(
          prev_key0_reg[106]), .Q(n3198));
   XNOR3X1 U5096 (.IN1(prev_key1_reg[106]), .IN2(new_sboxw[2]), .IN3(n3199), .Q(n2724));
   XNOR2X1 U5097 (.IN1(prev_key1_reg[42]), .IN2(prev_key1_reg[74]), .Q(n3199));
   AOI222X1 U5098 (.IN1(prev_key1_reg[42]), .IN2(n6949), .IN3(n7087), .IN4(key[42]), .IN5(
          key[170]), .IN6(n6703), .QN(n3196));
   AOI222X1 U5099 (.IN1(n2729), .IN2(n7053), .IN3(n2726), .IN4(n7143), .IN5(n2728), .IN6(
          n7101), .QN(n3201));
   XOR2X1 U5100 (.IN1(n3202), .IN2(n7615), .Q(n2728));
   XOR2X1 U5101 (.IN1(n3202), .IN2(n7613), .Q(n2726));
   XNOR3X1 U5102 (.IN1(prev_key0_reg[73]), .IN2(prev_key0_reg[41]), .IN3(
          prev_key0_reg[105]), .Q(n3202));
   XNOR3X1 U5103 (.IN1(prev_key1_reg[105]), .IN2(new_sboxw[1]), .IN3(n3203), .Q(n2729));
   XNOR2X1 U5104 (.IN1(prev_key1_reg[41]), .IN2(prev_key1_reg[73]), .Q(n3203));
   AOI222X1 U5105 (.IN1(prev_key1_reg[41]), .IN2(n6945), .IN3(n7087), .IN4(key[41]), .IN5(
          key[169]), .IN6(n6708), .QN(n3200));
   AOI222X1 U5106 (.IN1(n2734), .IN2(n7053), .IN3(n2731), .IN4(n7143), .IN5(n2733), .IN6(
          n7101), .QN(n3205));
   XOR2X1 U5107 (.IN1(n3206), .IN2(n7614), .Q(n2733));
   XOR2X1 U5108 (.IN1(n3206), .IN2(n7612), .Q(n2731));
   XNOR3X1 U5109 (.IN1(prev_key0_reg[72]), .IN2(prev_key0_reg[40]), .IN3(
          prev_key0_reg[104]), .Q(n3206));
   XNOR3X1 U5110 (.IN1(prev_key1_reg[104]), .IN2(new_sboxw[0]), .IN3(n3207), .Q(n2734));
   XNOR2X1 U5111 (.IN1(prev_key1_reg[40]), .IN2(prev_key1_reg[72]), .Q(n3207));
   AOI222X1 U5112 (.IN1(prev_key1_reg[40]), .IN2(n6948), .IN3(n7087), .IN4(key[40]), .IN5(
          key[168]), .IN6(n6707), .QN(n3204));
   AOI222X1 U5113 (.IN1(n2739), .IN2(n7053), .IN3(n2736), .IN4(n7143), .IN5(n2738), .IN6(
          n7101), .QN(n3209));
   XOR2X1 U5114 (.IN1(n3210), .IN2(n7598), .Q(n2738));
   XOR2X1 U5115 (.IN1(n3210), .IN2(n7621), .Q(n2736));
   XNOR3X1 U5116 (.IN1(prev_key0_reg[71]), .IN2(prev_key0_reg[39]), .IN3(
          prev_key0_reg[103]), .Q(n3210));
   XNOR3X1 U5117 (.IN1(prev_key1_reg[103]), .IN2(new_sboxw[31]), .IN3(n3211), .Q(n2739));
   XNOR2X1 U5118 (.IN1(prev_key1_reg[39]), .IN2(prev_key1_reg[71]), .Q(n3211));
   AOI222X1 U5119 (.IN1(prev_key1_reg[39]), .IN2(n6944), .IN3(n7087), .IN4(key[39]), .IN5(
          key[167]), .IN6(n6706), .QN(n3208));
   AOI222X1 U5120 (.IN1(n2744), .IN2(n7053), .IN3(n2741), .IN4(n7143), .IN5(n2743), .IN6(
          n7101), .QN(n3213));
   XOR2X1 U5121 (.IN1(n3214), .IN2(n7597), .Q(n2743));
   XOR2X1 U5122 (.IN1(n3214), .IN2(n7620), .Q(n2741));
   XNOR3X1 U5123 (.IN1(prev_key0_reg[70]), .IN2(prev_key0_reg[38]), .IN3(
          prev_key0_reg[102]), .Q(n3214));
   XNOR3X1 U5124 (.IN1(prev_key1_reg[102]), .IN2(new_sboxw[30]), .IN3(n3215), .Q(n2744));
   XNOR2X1 U5125 (.IN1(prev_key1_reg[38]), .IN2(prev_key1_reg[70]), .Q(n3215));
   AOI222X1 U5126 (.IN1(prev_key1_reg[38]), .IN2(n6945), .IN3(n7088), .IN4(key[38]), .IN5(
          key[166]), .IN6(n6705), .QN(n3212));
   AOI222X1 U5127 (.IN1(n2749), .IN2(n7053), .IN3(n2746), .IN4(n7143), .IN5(n2748), .IN6(
          n7101), .QN(n3217));
   XOR2X1 U5128 (.IN1(n3218), .IN2(n7596), .Q(n2748));
   XOR2X1 U5129 (.IN1(n3218), .IN2(n7619), .Q(n2746));
   XNOR3X1 U5130 (.IN1(prev_key0_reg[69]), .IN2(prev_key0_reg[37]), .IN3(
          prev_key0_reg[101]), .Q(n3218));
   XNOR3X1 U5131 (.IN1(prev_key1_reg[101]), .IN2(new_sboxw[29]), .IN3(n3219), .Q(n2749));
   XNOR2X1 U5132 (.IN1(prev_key1_reg[37]), .IN2(prev_key1_reg[69]), .Q(n3219));
   AOI222X1 U5133 (.IN1(prev_key1_reg[37]), .IN2(n6946), .IN3(n7088), .IN4(key[37]), .IN5(
          key[165]), .IN6(n6710), .QN(n3216));
   AOI222X1 U5134 (.IN1(n2754), .IN2(n7054), .IN3(n2751), .IN4(n7143), .IN5(n2753), .IN6(
          n7101), .QN(n3221));
   XOR2X1 U5135 (.IN1(n3222), .IN2(n7595), .Q(n2753));
   XOR2X1 U5136 (.IN1(n3222), .IN2(n7618), .Q(n2751));
   XNOR3X1 U5137 (.IN1(prev_key0_reg[68]), .IN2(prev_key0_reg[36]), .IN3(
          prev_key0_reg[100]), .Q(n3222));
   XNOR3X1 U5138 (.IN1(prev_key1_reg[100]), .IN2(new_sboxw[28]), .IN3(n3223), .Q(n2754));
   XNOR2X1 U5139 (.IN1(prev_key1_reg[36]), .IN2(prev_key1_reg[68]), .Q(n3223));
   AOI222X1 U5140 (.IN1(prev_key1_reg[36]), .IN2(n6945), .IN3(n7088), .IN4(key[36]), .IN5(
          key[164]), .IN6(n6709), .QN(n3220));
   AOI222X1 U5141 (.IN1(n2759), .IN2(n7054), .IN3(n2756), .IN4(n7143), .IN5(n2758), .IN6(
          n7100), .QN(n3225));
   XOR2X1 U5142 (.IN1(n3226), .IN2(n7594), .Q(n2758));
   XOR2X1 U5143 (.IN1(n3226), .IN2(n7617), .Q(n2756));
   XNOR3X1 U5144 (.IN1(prev_key0_reg[99]), .IN2(prev_key0_reg[67]), .IN3(prev_key0_reg[35])
          , .Q(n3226));
   XNOR3X1 U5145 (.IN1(prev_key1_reg[35]), .IN2(new_sboxw[27]), .IN3(n3227), .Q(n2759));
   XNOR2X1 U5146 (.IN1(prev_key1_reg[67]), .IN2(prev_key1_reg[99]), .Q(n3227));
   AOI222X1 U5147 (.IN1(prev_key1_reg[35]), .IN2(n6946), .IN3(n7088), .IN4(key[35]), .IN5(
          key[163]), .IN6(n6704), .QN(n3224));
   AOI222X1 U5148 (.IN1(n2764), .IN2(n7054), .IN3(n2761), .IN4(n7143), .IN5(n2763), .IN6(
          n7100), .QN(n3229));
   XOR2X1 U5149 (.IN1(n3230), .IN2(n7593), .Q(n2763));
   XOR2X1 U5150 (.IN1(n3230), .IN2(n7616), .Q(n2761));
   XNOR3X1 U5151 (.IN1(prev_key0_reg[98]), .IN2(prev_key0_reg[66]), .IN3(prev_key0_reg[34])
          , .Q(n3230));
   XNOR3X1 U5152 (.IN1(prev_key1_reg[34]), .IN2(new_sboxw[26]), .IN3(n3231), .Q(n2764));
   XNOR2X1 U5153 (.IN1(prev_key1_reg[66]), .IN2(prev_key1_reg[98]), .Q(n3231));
   AOI222X1 U5154 (.IN1(prev_key1_reg[34]), .IN2(n6947), .IN3(n7088), .IN4(key[34]), .IN5(
          key[162]), .IN6(n6703), .QN(n3228));
   AOI222X1 U5155 (.IN1(n2769), .IN2(n7054), .IN3(n2766), .IN4(n7143), .IN5(n2768), .IN6(
          n7100), .QN(n3233));
   XOR2X1 U5156 (.IN1(n3234), .IN2(n7592), .Q(n2768));
   XOR2X1 U5157 (.IN1(n3234), .IN2(n7615), .Q(n2766));
   XNOR3X1 U5158 (.IN1(prev_key0_reg[97]), .IN2(prev_key0_reg[65]), .IN3(prev_key0_reg[33])
          , .Q(n3234));
   XNOR3X1 U5159 (.IN1(prev_key1_reg[33]), .IN2(new_sboxw[25]), .IN3(n3235), .Q(n2769));
   XNOR2X1 U5160 (.IN1(prev_key1_reg[65]), .IN2(prev_key1_reg[97]), .Q(n3235));
   AOI222X1 U5161 (.IN1(prev_key1_reg[33]), .IN2(n6948), .IN3(n7088), .IN4(key[33]), .IN5(
          key[161]), .IN6(n6711), .QN(n3232));
   AOI222X1 U5162 (.IN1(n2774), .IN2(n7054), .IN3(n2771), .IN4(n7143), .IN5(n2773), .IN6(
          n7100), .QN(n3237));
   XOR2X1 U5163 (.IN1(n3238), .IN2(n7591), .Q(n2773));
   XOR2X1 U5164 (.IN1(n3238), .IN2(n7614), .Q(n2771));
   XNOR3X1 U5165 (.IN1(prev_key0_reg[96]), .IN2(prev_key0_reg[64]), .IN3(prev_key0_reg[32])
          , .Q(n3238));
   XNOR3X1 U5166 (.IN1(prev_key1_reg[32]), .IN2(new_sboxw[24]), .IN3(n3239), .Q(n2774));
   XNOR2X1 U5167 (.IN1(prev_key1_reg[64]), .IN2(prev_key1_reg[96]), .Q(n3239));
   AOI222X1 U5168 (.IN1(prev_key1_reg[32]), .IN2(n6949), .IN3(n7088), .IN4(key[32]), .IN5(
          key[160]), .IN6(n6710), .QN(n3236));
   AOI222X1 U5169 (.IN1(n2779), .IN2(n7054), .IN3(n2776), .IN4(n7144), .IN5(n2778), .IN6(
          n7100), .QN(n3241));
   XOR2X1 U5170 (.IN1(n3242), .IN2(n7590), .Q(n2778));
   XOR2X1 U5171 (.IN1(n3242), .IN2(n7598), .Q(n2776));
   XNOR3X1 U5172 (.IN1(prev_key0_reg[31]), .IN2(n2215), .IN3(n3243), .Q(n3242));
   XNOR2X1 U5173 (.IN1(prev_key0_reg[63]), .IN2(prev_key0_reg[95]), .Q(n3243));
   XNOR3X1 U5174 (.IN1(prev_key1_reg[127]), .IN2(n3018), .IN3(n3244), .Q(n2779));
   XNOR3X1 U5175 (.IN1(sboxw[31]), .IN2(prev_key1_reg[95]), .IN3(prev_key1_reg[63]), .Q(
          n3244));
   XOR2X1 U5176 (.IN1(new_sboxw[23]), .IN2(rcon_reg[7]), .Q(n3018));
   AOI222X1 U5177 (.IN1(sboxw[31]), .IN2(n6947), .IN3(n7088), .IN4(key[31]), .IN5(key[159])
          , .IN6(n6710), .QN(n3240));
   AOI222X1 U5178 (.IN1(n2784), .IN2(n7054), .IN3(n2781), .IN4(n7144), .IN5(n2783), .IN6(
          n7100), .QN(n3246));
   XOR2X1 U5179 (.IN1(n3247), .IN2(n2948), .Q(n2783));
   XOR2X1 U5180 (.IN1(n3247), .IN2(n7597), .Q(n2781));
   XNOR3X1 U5181 (.IN1(prev_key0_reg[30]), .IN2(n2216), .IN3(n3248), .Q(n3247));
   XNOR2X1 U5182 (.IN1(prev_key0_reg[62]), .IN2(prev_key0_reg[94]), .Q(n3248));
   XNOR3X1 U5183 (.IN1(prev_key1_reg[126]), .IN2(n7589), .IN3(n3249), .Q(n2784));
   XNOR3X1 U5184 (.IN1(sboxw[30]), .IN2(prev_key1_reg[94]), .IN3(prev_key1_reg[62]), .Q(
          n3249));
   XOR2X1 U5185 (.IN1(rcon_reg[6]), .IN2(n7605), .Q(n2948));
   AOI222X1 U5186 (.IN1(sboxw[30]), .IN2(n6950), .IN3(n7088), .IN4(key[30]), .IN5(key[158])
          , .IN6(n6709), .QN(n3245));
   AOI222X1 U5187 (.IN1(n2789), .IN2(n7054), .IN3(n2786), .IN4(n7144), .IN5(n2788), .IN6(
          n7100), .QN(n3251));
   XOR2X1 U5188 (.IN1(n3252), .IN2(n2951), .Q(n2788));
   XOR2X1 U5189 (.IN1(n3252), .IN2(n7596), .Q(n2786));
   XNOR3X1 U5190 (.IN1(prev_key0_reg[29]), .IN2(n2217), .IN3(n3253), .Q(n3252));
   XNOR2X1 U5191 (.IN1(prev_key0_reg[61]), .IN2(prev_key0_reg[93]), .Q(n3253));
   XNOR3X1 U5192 (.IN1(prev_key1_reg[125]), .IN2(n7588), .IN3(n3254), .Q(n2789));
   XNOR3X1 U5193 (.IN1(sboxw[29]), .IN2(prev_key1_reg[93]), .IN3(prev_key1_reg[61]), .Q(
          n3254));
   XOR2X1 U5194 (.IN1(rcon_reg[5]), .IN2(n7604), .Q(n2951));
   AOI222X1 U5195 (.IN1(sboxw[29]), .IN2(n6951), .IN3(n7088), .IN4(key[29]), .IN5(key[157])
          , .IN6(n6708), .QN(n3250));
   AOI222X1 U5196 (.IN1(n2794), .IN2(n7054), .IN3(n2791), .IN4(n7144), .IN5(n2793), .IN6(
          n7100), .QN(n3256));
   XOR2X1 U5197 (.IN1(n3257), .IN2(n2954), .Q(n2793));
   XOR2X1 U5198 (.IN1(n3257), .IN2(n7595), .Q(n2791));
   XNOR3X1 U5199 (.IN1(prev_key0_reg[28]), .IN2(n2218), .IN3(n3258), .Q(n3257));
   XNOR2X1 U5200 (.IN1(prev_key0_reg[60]), .IN2(prev_key0_reg[92]), .Q(n3258));
   XNOR3X1 U5201 (.IN1(prev_key1_reg[124]), .IN2(n7587), .IN3(n3259), .Q(n2794));
   XNOR3X1 U5202 (.IN1(sboxw[28]), .IN2(prev_key1_reg[92]), .IN3(prev_key1_reg[60]), .Q(
          n3259));
   XOR2X1 U5203 (.IN1(rcon_reg[4]), .IN2(n7603), .Q(n2954));
   AOI222X1 U5204 (.IN1(sboxw[28]), .IN2(n6952), .IN3(n7088), .IN4(key[28]), .IN5(key[156])
          , .IN6(n6707), .QN(n3255));
   AOI222X1 U5205 (.IN1(n2799), .IN2(n7054), .IN3(n2796), .IN4(n7144), .IN5(n2798), .IN6(
          n7100), .QN(n3261));
   XOR2X1 U5206 (.IN1(n3262), .IN2(n2957), .Q(n2798));
   XOR2X1 U5207 (.IN1(n3262), .IN2(n7594), .Q(n2796));
   XNOR3X1 U5208 (.IN1(prev_key0_reg[27]), .IN2(n2219), .IN3(n3263), .Q(n3262));
   XNOR2X1 U5209 (.IN1(prev_key0_reg[59]), .IN2(prev_key0_reg[91]), .Q(n3263));
   XNOR3X1 U5210 (.IN1(prev_key1_reg[123]), .IN2(n7586), .IN3(n3264), .Q(n2799));
   XNOR3X1 U5211 (.IN1(sboxw[27]), .IN2(prev_key1_reg[91]), .IN3(prev_key1_reg[59]), .Q(
          n3264));
   XOR2X1 U5212 (.IN1(rcon_reg[3]), .IN2(n7602), .Q(n2957));
   AOI222X1 U5213 (.IN1(sboxw[27]), .IN2(n6953), .IN3(n7088), .IN4(key[27]), .IN5(key[155])
          , .IN6(n6708), .QN(n3260));
   AOI222X1 U5214 (.IN1(n2804), .IN2(n7054), .IN3(n2801), .IN4(n7144), .IN5(n2803), .IN6(
          n7100), .QN(n3266));
   XOR2X1 U5215 (.IN1(n3267), .IN2(n2960), .Q(n2803));
   XOR2X1 U5216 (.IN1(n3267), .IN2(n7593), .Q(n2801));
   XNOR3X1 U5217 (.IN1(prev_key0_reg[26]), .IN2(n2220), .IN3(n3268), .Q(n3267));
   XNOR2X1 U5218 (.IN1(prev_key0_reg[58]), .IN2(prev_key0_reg[90]), .Q(n3268));
   XNOR3X1 U5219 (.IN1(prev_key1_reg[122]), .IN2(n7585), .IN3(n3269), .Q(n2804));
   XNOR3X1 U5220 (.IN1(sboxw[26]), .IN2(prev_key1_reg[90]), .IN3(prev_key1_reg[58]), .Q(
          n3269));
   XOR2X1 U5221 (.IN1(rcon_reg[2]), .IN2(n7601), .Q(n2960));
   AOI222X1 U5222 (.IN1(sboxw[26]), .IN2(n6954), .IN3(n7088), .IN4(key[26]), .IN5(key[154])
          , .IN6(n6707), .QN(n3265));
   AOI222X1 U5223 (.IN1(n2809), .IN2(n7054), .IN3(n2806), .IN4(n7144), .IN5(n2808), .IN6(
          n7100), .QN(n3271));
   XOR2X1 U5224 (.IN1(n3272), .IN2(n2963), .Q(n2808));
   XOR2X1 U5225 (.IN1(n3272), .IN2(n7592), .Q(n2806));
   XNOR3X1 U5226 (.IN1(prev_key0_reg[25]), .IN2(n2221), .IN3(n3273), .Q(n3272));
   XNOR2X1 U5227 (.IN1(prev_key0_reg[57]), .IN2(prev_key0_reg[89]), .Q(n3273));
   XNOR3X1 U5228 (.IN1(prev_key1_reg[121]), .IN2(n7584), .IN3(n3274), .Q(n2809));
   XNOR3X1 U5229 (.IN1(sboxw[25]), .IN2(prev_key1_reg[89]), .IN3(prev_key1_reg[57]), .Q(
          n3274));
   XOR2X1 U5230 (.IN1(rcon_reg[1]), .IN2(n7600), .Q(n2963));
   AOI222X1 U5231 (.IN1(sboxw[25]), .IN2(n6948), .IN3(n7088), .IN4(key[25]), .IN5(key[153])
          , .IN6(n6706), .QN(n3270));
   AOI222X1 U5232 (.IN1(n2814), .IN2(n7054), .IN3(n2811), .IN4(n7144), .IN5(n2813), .IN6(
          n7100), .QN(n3276));
   XOR2X1 U5233 (.IN1(n3277), .IN2(n2966), .Q(n2813));
   XOR2X1 U5234 (.IN1(n3277), .IN2(n7591), .Q(n2811));
   XNOR3X1 U5235 (.IN1(prev_key0_reg[24]), .IN2(n2222), .IN3(n3278), .Q(n3277));
   XNOR2X1 U5236 (.IN1(prev_key0_reg[56]), .IN2(prev_key0_reg[88]), .Q(n3278));
   XOR2X1 U5239 (.IN1(rcon_reg[0]), .IN2(n7599), .Q(n2966));
   AOI222X1 U5240 (.IN1(sboxw[24]), .IN2(n6945), .IN3(n7089), .IN4(key[24]), .IN5(key[152])
          , .IN6(n6705), .QN(n3275));
   AOI222X1 U5241 (.IN1(n2819), .IN2(n7054), .IN3(n2816), .IN4(n7144), .IN5(n2818), .IN6(
          n7099), .QN(n3281));
   XOR2X1 U5242 (.IN1(n3282), .IN2(n7611), .Q(n2818));
   XNOR2X1 U5243 (.IN1(n3282), .IN2(new_sboxw[23]), .Q(n2816));
   XNOR3X1 U5244 (.IN1(prev_key0_reg[23]), .IN2(n2223), .IN3(n3283), .Q(n3282));
   XNOR2X1 U5245 (.IN1(prev_key0_reg[55]), .IN2(prev_key0_reg[87]), .Q(n3283));
   XNOR3X1 U5246 (.IN1(prev_key1_reg[119]), .IN2(new_sboxw[15]), .IN3(n3284), .Q(n2819));
   XNOR3X1 U5247 (.IN1(sboxw[23]), .IN2(prev_key1_reg[87]), .IN3(prev_key1_reg[55]), .Q(
          n3284));
   AOI222X1 U5248 (.IN1(sboxw[23]), .IN2(n6954), .IN3(n7089), .IN4(key[23]), .IN5(key[151])
          , .IN6(n6704), .QN(n3280));
   AOI222X1 U5249 (.IN1(n2824), .IN2(n7054), .IN3(n2821), .IN4(n7144), .IN5(n2823), .IN6(
          n7099), .QN(n3286));
   XOR2X1 U5250 (.IN1(n3287), .IN2(n6701), .Q(n2823));
   XOR2X1 U5251 (.IN1(n3287), .IN2(n7605), .Q(n2821));
   XNOR3X1 U5252 (.IN1(prev_key0_reg[22]), .IN2(n2224), .IN3(n3288), .Q(n3287));
   XNOR2X1 U5253 (.IN1(prev_key0_reg[54]), .IN2(prev_key0_reg[86]), .Q(n3288));
   XNOR3X1 U5254 (.IN1(prev_key1_reg[118]), .IN2(new_sboxw[14]), .IN3(n3289), .Q(n2824));
   XNOR3X1 U5255 (.IN1(sboxw[22]), .IN2(prev_key1_reg[86]), .IN3(prev_key1_reg[54]), .Q(
          n3289));
   AOI222X1 U5256 (.IN1(sboxw[22]), .IN2(n6944), .IN3(n7089), .IN4(key[22]), .IN5(key[150])
          , .IN6(n6703), .QN(n3285));
   AOI222X1 U5257 (.IN1(n2829), .IN2(n7054), .IN3(n2826), .IN4(n7144), .IN5(n2828), .IN6(
          n7099), .QN(n3291));
   XOR2X1 U5258 (.IN1(n3292), .IN2(n7609), .Q(n2828));
   XOR2X1 U5259 (.IN1(n3292), .IN2(n7604), .Q(n2826));
   XNOR3X1 U5260 (.IN1(prev_key0_reg[21]), .IN2(n2225), .IN3(n3293), .Q(n3292));
   XNOR2X1 U5261 (.IN1(prev_key0_reg[53]), .IN2(prev_key0_reg[85]), .Q(n3293));
   XNOR3X1 U5262 (.IN1(prev_key1_reg[117]), .IN2(new_sboxw[13]), .IN3(n3294), .Q(n2829));
   XNOR3X1 U5263 (.IN1(sboxw[21]), .IN2(prev_key1_reg[85]), .IN3(prev_key1_reg[53]), .Q(
          n3294));
   AOI222X1 U5264 (.IN1(sboxw[21]), .IN2(n6947), .IN3(n7089), .IN4(key[21]), .IN5(key[149])
          , .IN6(n6711), .QN(n3290));
   AOI222X1 U5265 (.IN1(n2834), .IN2(n7054), .IN3(n2831), .IN4(n7144), .IN5(n2833), .IN6(
          n7099), .QN(n3296));
   XOR2X1 U5266 (.IN1(n3297), .IN2(n7608), .Q(n2833));
   XOR2X1 U5267 (.IN1(n3297), .IN2(n7603), .Q(n2831));
   XNOR3X1 U5268 (.IN1(prev_key0_reg[20]), .IN2(n2226), .IN3(n3298), .Q(n3297));
   XNOR2X1 U5269 (.IN1(prev_key0_reg[52]), .IN2(prev_key0_reg[84]), .Q(n3298));
   XNOR3X1 U5270 (.IN1(prev_key1_reg[116]), .IN2(new_sboxw[12]), .IN3(n3299), .Q(n2834));
   XNOR3X1 U5271 (.IN1(sboxw[20]), .IN2(prev_key1_reg[84]), .IN3(prev_key1_reg[52]), .Q(
          n3299));
   AOI222X1 U5272 (.IN1(sboxw[20]), .IN2(n6948), .IN3(n7089), .IN4(key[20]), .IN5(key[148])
          , .IN6(n2945), .QN(n3295));
   AOI222X1 U5273 (.IN1(n2839), .IN2(n7055), .IN3(n2836), .IN4(n7144), .IN5(n2838), .IN6(
          n7099), .QN(n3301));
   XOR2X1 U5274 (.IN1(n3302), .IN2(n7607), .Q(n2838));
   XOR2X1 U5275 (.IN1(n3302), .IN2(n7602), .Q(n2836));
   XNOR3X1 U5276 (.IN1(prev_key0_reg[19]), .IN2(n2227), .IN3(n3303), .Q(n3302));
   XNOR2X1 U5277 (.IN1(prev_key0_reg[51]), .IN2(prev_key0_reg[83]), .Q(n3303));
   XNOR3X1 U5278 (.IN1(prev_key1_reg[115]), .IN2(new_sboxw[11]), .IN3(n3304), .Q(n2839));
   XNOR3X1 U5279 (.IN1(sboxw[19]), .IN2(prev_key1_reg[83]), .IN3(prev_key1_reg[51]), .Q(
          n3304));
   AOI222X1 U5280 (.IN1(sboxw[19]), .IN2(n6949), .IN3(n7089), .IN4(key[19]), .IN5(key[147])
          , .IN6(n6710), .QN(n3300));
   AOI222X1 U5281 (.IN1(n2844), .IN2(n7055), .IN3(n2841), .IN4(n7145), .IN5(n2843), .IN6(
          n7099), .QN(n3306));
   XOR2X1 U5282 (.IN1(n3307), .IN2(n7606), .Q(n2843));
   XOR2X1 U5283 (.IN1(n3307), .IN2(n7601), .Q(n2841));
   XNOR3X1 U5284 (.IN1(prev_key0_reg[18]), .IN2(n2228), .IN3(n3308), .Q(n3307));
   XNOR2X1 U5285 (.IN1(prev_key0_reg[50]), .IN2(prev_key0_reg[82]), .Q(n3308));
   XNOR3X1 U5286 (.IN1(prev_key1_reg[114]), .IN2(new_sboxw[10]), .IN3(n3309), .Q(n2844));
   XNOR3X1 U5287 (.IN1(sboxw[18]), .IN2(prev_key1_reg[82]), .IN3(prev_key1_reg[50]), .Q(
          n3309));
   AOI222X1 U5288 (.IN1(sboxw[18]), .IN2(n6946), .IN3(n7089), .IN4(key[18]), .IN5(key[146])
          , .IN6(n6709), .QN(n3305));
   AOI222X1 U5289 (.IN1(n2849), .IN2(n7055), .IN3(n2846), .IN4(n7145), .IN5(n2848), .IN6(
          n7099), .QN(n3311));
   XOR2X1 U5290 (.IN1(n3312), .IN2(n7613), .Q(n2848));
   XOR2X1 U5291 (.IN1(n3312), .IN2(n7600), .Q(n2846));
   XNOR3X1 U5292 (.IN1(prev_key0_reg[17]), .IN2(n2229), .IN3(n3313), .Q(n3312));
   XNOR2X1 U5293 (.IN1(prev_key0_reg[49]), .IN2(prev_key0_reg[81]), .Q(n3313));
   XNOR3X1 U5294 (.IN1(prev_key1_reg[113]), .IN2(new_sboxw[9]), .IN3(n3314), .Q(n2849));
   XNOR3X1 U5295 (.IN1(sboxw[17]), .IN2(prev_key1_reg[81]), .IN3(prev_key1_reg[49]), .Q(
          n3314));
   AOI222X1 U5296 (.IN1(sboxw[17]), .IN2(n6955), .IN3(n7089), .IN4(key[17]), .IN5(key[145])
          , .IN6(n6706), .QN(n3310));
   AOI222X1 U5297 (.IN1(n2854), .IN2(n7055), .IN3(n2851), .IN4(n7145), .IN5(n2853), .IN6(
          n7099), .QN(n3316));
   XOR2X1 U5298 (.IN1(n3317), .IN2(n7612), .Q(n2853));
   XOR2X1 U5299 (.IN1(n3317), .IN2(n7599), .Q(n2851));
   XNOR3X1 U5300 (.IN1(prev_key0_reg[16]), .IN2(n2230), .IN3(n3318), .Q(n3317));
   XNOR2X1 U5301 (.IN1(prev_key0_reg[48]), .IN2(prev_key0_reg[80]), .Q(n3318));
   XNOR3X1 U5302 (.IN1(prev_key1_reg[112]), .IN2(new_sboxw[8]), .IN3(n3319), .Q(n2854));
   XNOR3X1 U5303 (.IN1(sboxw[16]), .IN2(prev_key1_reg[80]), .IN3(prev_key1_reg[48]), .Q(
          n3319));
   AOI222X1 U5304 (.IN1(sboxw[16]), .IN2(n6946), .IN3(n7089), .IN4(key[16]), .IN5(key[144])
          , .IN6(n6705), .QN(n3315));
   AOI222X1 U5305 (.IN1(n2859), .IN2(n7055), .IN3(n2856), .IN4(n7145), .IN5(n2858), .IN6(
          n7099), .QN(n3321));
   XOR2X1 U5306 (.IN1(n3322), .IN2(n7621), .Q(n2858));
   XOR2X1 U5307 (.IN1(n3322), .IN2(n7611), .Q(n2856));
   XOR3X1 U5308 (.IN1(prev_key0_reg[15]), .IN2(prev_key0_reg[111]), .IN3(n3323), .Q(n3322)
          );
   XNOR2X1 U5309 (.IN1(prev_key0_reg[47]), .IN2(prev_key0_reg[79]), .Q(n3323));
   AOI222X1 U5312 (.IN1(sboxw[15]), .IN2(n6955), .IN3(n7089), .IN4(key[15]), .IN5(key[143])
          , .IN6(n6708), .QN(n3320));
   AOI222X1 U5313 (.IN1(n2864), .IN2(n7055), .IN3(n2861), .IN4(n7145), .IN5(n2863), .IN6(
          n7099), .QN(n3326));
   XOR2X1 U5314 (.IN1(n3327), .IN2(n7620), .Q(n2863));
   XOR2X1 U5315 (.IN1(n3327), .IN2(n6701), .Q(n2861));
   XOR3X1 U5316 (.IN1(prev_key0_reg[14]), .IN2(prev_key0_reg[110]), .IN3(n3328), .Q(n3327)
          );
   XNOR2X1 U5317 (.IN1(prev_key0_reg[46]), .IN2(prev_key0_reg[78]), .Q(n3328));
   XNOR3X1 U5318 (.IN1(prev_key1_reg[110]), .IN2(new_sboxw[6]), .IN3(n3329), .Q(n2864));
   XNOR3X1 U5319 (.IN1(sboxw[14]), .IN2(prev_key1_reg[78]), .IN3(prev_key1_reg[46]), .Q(
          n3329));
   AOI222X1 U5320 (.IN1(sboxw[14]), .IN2(n6949), .IN3(n7089), .IN4(key[14]), .IN5(key[142])
          , .IN6(n6707), .QN(n3325));
   AOI222X1 U5321 (.IN1(n2869), .IN2(n7055), .IN3(n2866), .IN4(n7145), .IN5(n2868), .IN6(
          n7099), .QN(n3331));
   XOR2X1 U5322 (.IN1(n3332), .IN2(n7619), .Q(n2868));
   XOR2X1 U5323 (.IN1(n3332), .IN2(n7609), .Q(n2866));
   XOR3X1 U5324 (.IN1(prev_key0_reg[13]), .IN2(prev_key0_reg[109]), .IN3(n3333), .Q(n3332)
          );
   XNOR2X1 U5325 (.IN1(prev_key0_reg[45]), .IN2(prev_key0_reg[77]), .Q(n3333));
   AOI222X1 U5328 (.IN1(sboxw[13]), .IN2(n6944), .IN3(n7089), .IN4(key[13]), .IN5(key[141])
          , .IN6(n6706), .QN(n3330));
   AOI222X1 U5329 (.IN1(n2874), .IN2(n7055), .IN3(n2871), .IN4(n7145), .IN5(n2873), .IN6(
          n7099), .QN(n3336));
   XOR2X1 U5330 (.IN1(n3337), .IN2(n7618), .Q(n2873));
   XOR2X1 U5331 (.IN1(n3337), .IN2(n7608), .Q(n2871));
   XOR3X1 U5332 (.IN1(prev_key0_reg[12]), .IN2(prev_key0_reg[108]), .IN3(n3338), .Q(n3337)
          );
   XNOR2X1 U5333 (.IN1(prev_key0_reg[44]), .IN2(prev_key0_reg[76]), .Q(n3338));
   XNOR3X1 U5334 (.IN1(prev_key1_reg[108]), .IN2(new_sboxw[4]), .IN3(n3339), .Q(n2874));
   XNOR3X1 U5335 (.IN1(sboxw[12]), .IN2(prev_key1_reg[76]), .IN3(prev_key1_reg[44]), .Q(
          n3339));
   AOI222X1 U5336 (.IN1(sboxw[12]), .IN2(n6945), .IN3(n7089), .IN4(key[12]), .IN5(key[140])
          , .IN6(n6705), .QN(n3335));
   AOI222X1 U5337 (.IN1(n2879), .IN2(n7055), .IN3(n2876), .IN4(n7145), .IN5(n2878), .IN6(
          n7098), .QN(n3341));
   XOR2X1 U5338 (.IN1(n3342), .IN2(n7617), .Q(n2878));
   XOR2X1 U5339 (.IN1(n3342), .IN2(n7607), .Q(n2876));
   XOR3X1 U5340 (.IN1(prev_key0_reg[11]), .IN2(prev_key0_reg[107]), .IN3(n3343), .Q(n3342)
          );
   XNOR2X1 U5341 (.IN1(prev_key0_reg[43]), .IN2(prev_key0_reg[75]), .Q(n3343));
   XNOR3X1 U5342 (.IN1(prev_key1_reg[107]), .IN2(new_sboxw[3]), .IN3(n3344), .Q(n2879));
   XNOR3X1 U5343 (.IN1(sboxw[11]), .IN2(prev_key1_reg[75]), .IN3(prev_key1_reg[43]), .Q(
          n3344));
   AOI222X1 U5344 (.IN1(sboxw[11]), .IN2(n6946), .IN3(n7089), .IN4(key[11]), .IN5(key[139])
          , .IN6(n6704), .QN(n3340));
   AOI222X1 U5345 (.IN1(n2884), .IN2(n7055), .IN3(n2881), .IN4(n7145), .IN5(n2883), .IN6(
          n7098), .QN(n3346));
   XOR2X1 U5346 (.IN1(n3347), .IN2(n7616), .Q(n2883));
   XOR2X1 U5347 (.IN1(n3347), .IN2(n7606), .Q(n2881));
   XOR3X1 U5348 (.IN1(prev_key0_reg[10]), .IN2(prev_key0_reg[106]), .IN3(n3348), .Q(n3347)
          );
   XNOR2X1 U5349 (.IN1(prev_key0_reg[42]), .IN2(prev_key0_reg[74]), .Q(n3348));
   AOI222X1 U5352 (.IN1(sboxw[10]), .IN2(n6947), .IN3(n7090), .IN4(key[10]), .IN5(key[138])
          , .IN6(n6703), .QN(n3345));
   AOI222X1 U5353 (.IN1(n2889), .IN2(n7055), .IN3(n2886), .IN4(n7145), .IN5(n2888), .IN6(
          n7098), .QN(n3351));
   XOR2X1 U5354 (.IN1(n3352), .IN2(n7615), .Q(n2888));
   XOR2X1 U5355 (.IN1(n3352), .IN2(n7613), .Q(n2886));
   XOR3X1 U5356 (.IN1(prev_key0_reg[41]), .IN2(prev_key0_reg[105]), .IN3(n3353), .Q(n3352)
          );
   XNOR2X1 U5357 (.IN1(prev_key0_reg[9]), .IN2(prev_key0_reg[73]), .Q(n3353));
   XNOR3X1 U5358 (.IN1(prev_key1_reg[105]), .IN2(new_sboxw[1]), .IN3(n3354), .Q(n2889));
   XNOR3X1 U5359 (.IN1(sboxw[9]), .IN2(prev_key1_reg[73]), .IN3(prev_key1_reg[41]), .Q(
          n3354));
   AOI222X1 U5360 (.IN1(sboxw[9]), .IN2(n6948), .IN3(n7090), .IN4(key[9]), .IN5(key[137])
          , .IN6(n6711), .QN(n3350));
   AOI222X1 U5361 (.IN1(n2894), .IN2(n7055), .IN3(n2891), .IN4(n7145), .IN5(n2893), .IN6(
          n7098), .QN(n3356));
   XOR2X1 U5362 (.IN1(n3357), .IN2(n7614), .Q(n2893));
   XOR2X1 U5363 (.IN1(n3357), .IN2(n7612), .Q(n2891));
   XOR3X1 U5364 (.IN1(prev_key0_reg[40]), .IN2(prev_key0_reg[104]), .IN3(n3358), .Q(n3357)
          );
   XNOR2X1 U5365 (.IN1(prev_key0_reg[8]), .IN2(prev_key0_reg[72]), .Q(n3358));
   XNOR3X1 U5366 (.IN1(prev_key1_reg[104]), .IN2(new_sboxw[0]), .IN3(n3359), .Q(n2894));
   XNOR3X1 U5367 (.IN1(sboxw[8]), .IN2(prev_key1_reg[72]), .IN3(prev_key1_reg[40]), .Q(
          n3359));
   AOI222X1 U5368 (.IN1(sboxw[8]), .IN2(n6949), .IN3(n7090), .IN4(key[8]), .IN5(key[136])
          , .IN6(n2945), .QN(n3355));
   AOI222X1 U5369 (.IN1(n2899), .IN2(n7055), .IN3(n2896), .IN4(n7145), .IN5(n2898), .IN6(
          n7098), .QN(n3361));
   XOR2X1 U5370 (.IN1(n3362), .IN2(n7598), .Q(n2898));
   XOR2X1 U5371 (.IN1(n3362), .IN2(n7621), .Q(n2896));
   XOR3X1 U5372 (.IN1(prev_key0_reg[39]), .IN2(prev_key0_reg[103]), .IN3(n3363), .Q(n3362)
          );
   XNOR2X1 U5373 (.IN1(prev_key0_reg[7]), .IN2(prev_key0_reg[71]), .Q(n3363));
   XNOR3X1 U5374 (.IN1(prev_key1_reg[103]), .IN2(new_sboxw[31]), .IN3(n3364), .Q(n2899));
   XNOR3X1 U5375 (.IN1(sboxw[7]), .IN2(prev_key1_reg[71]), .IN3(prev_key1_reg[39]), .Q(
          n3364));
   AOI222X1 U5376 (.IN1(sboxw[7]), .IN2(n6948), .IN3(n7090), .IN4(key[7]), .IN5(key[135])
          , .IN6(n6706), .QN(n3360));
   AOI222X1 U5377 (.IN1(n2904), .IN2(n7055), .IN3(n2901), .IN4(n7145), .IN5(n2903), .IN6(
          n7098), .QN(n3366));
   XOR2X1 U5378 (.IN1(n3367), .IN2(n7597), .Q(n2903));
   XOR2X1 U5379 (.IN1(n3367), .IN2(n7620), .Q(n2901));
   XOR3X1 U5380 (.IN1(prev_key0_reg[38]), .IN2(prev_key0_reg[102]), .IN3(n3368), .Q(n3367)
          );
   XNOR2X1 U5381 (.IN1(prev_key0_reg[6]), .IN2(prev_key0_reg[70]), .Q(n3368));
   XNOR3X1 U5382 (.IN1(prev_key1_reg[102]), .IN2(new_sboxw[30]), .IN3(n3369), .Q(n2904));
   XNOR3X1 U5383 (.IN1(sboxw[6]), .IN2(prev_key1_reg[70]), .IN3(prev_key1_reg[38]), .Q(
          n3369));
   AOI222X1 U5384 (.IN1(sboxw[6]), .IN2(n6955), .IN3(n7090), .IN4(key[6]), .IN5(key[134])
          , .IN6(n6705), .QN(n3365));
   AOI222X1 U5385 (.IN1(n2909), .IN2(n7055), .IN3(n2906), .IN4(n7146), .IN5(n2908), .IN6(
          n7098), .QN(n3371));
   XOR2X1 U5386 (.IN1(n3372), .IN2(n7596), .Q(n2908));
   XOR2X1 U5387 (.IN1(n3372), .IN2(n7619), .Q(n2906));
   XOR3X1 U5388 (.IN1(prev_key0_reg[37]), .IN2(prev_key0_reg[101]), .IN3(n3373), .Q(n3372)
          );
   XNOR2X1 U5389 (.IN1(prev_key0_reg[5]), .IN2(prev_key0_reg[69]), .Q(n3373));
   XNOR3X1 U5390 (.IN1(prev_key1_reg[101]), .IN2(new_sboxw[29]), .IN3(n3374), .Q(n2909));
   XNOR3X1 U5391 (.IN1(sboxw[5]), .IN2(prev_key1_reg[69]), .IN3(prev_key1_reg[37]), .Q(
          n3374));
   AOI222X1 U5392 (.IN1(sboxw[5]), .IN2(n6945), .IN3(n7090), .IN4(key[5]), .IN5(key[133])
          , .IN6(n6704), .QN(n3370));
   AOI222X1 U5393 (.IN1(n2914), .IN2(n7055), .IN3(n2911), .IN4(n7146), .IN5(n2913), .IN6(
          n7098), .QN(n3376));
   XOR2X1 U5394 (.IN1(n3377), .IN2(n7595), .Q(n2913));
   XOR2X1 U5395 (.IN1(n3377), .IN2(n7618), .Q(n2911));
   XOR3X1 U5396 (.IN1(prev_key0_reg[36]), .IN2(prev_key0_reg[100]), .IN3(n3378), .Q(n3377)
          );
   XNOR2X1 U5397 (.IN1(prev_key0_reg[4]), .IN2(prev_key0_reg[68]), .Q(n3378));
   XNOR3X1 U5398 (.IN1(prev_key1_reg[100]), .IN2(new_sboxw[28]), .IN3(n3379), .Q(n2914));
   XNOR3X1 U5399 (.IN1(sboxw[4]), .IN2(prev_key1_reg[68]), .IN3(prev_key1_reg[36]), .Q(
          n3379));
   AOI222X1 U5400 (.IN1(sboxw[4]), .IN2(n6946), .IN3(n7090), .IN4(key[4]), .IN5(key[132])
          , .IN6(n6703), .QN(n3375));
   AOI222X1 U5401 (.IN1(n2919), .IN2(n7055), .IN3(n2916), .IN4(n7146), .IN5(n2918), .IN6(
          n7098), .QN(n3381));
   XOR2X1 U5402 (.IN1(n3382), .IN2(n7594), .Q(n2918));
   XOR2X1 U5403 (.IN1(n3382), .IN2(n7617), .Q(n2916));
   XOR3X1 U5404 (.IN1(prev_key0_reg[99]), .IN2(prev_key0_reg[67]), .IN3(n3383), .Q(n3382)
          );
   XNOR2X1 U5405 (.IN1(prev_key0_reg[35]), .IN2(prev_key0_reg[3]), .Q(n3383));
   XNOR3X1 U5406 (.IN1(prev_key1_reg[35]), .IN2(new_sboxw[27]), .IN3(n3384), .Q(n2919));
   XNOR3X1 U5407 (.IN1(sboxw[3]), .IN2(prev_key1_reg[99]), .IN3(prev_key1_reg[67]), .Q(
          n3384));
   AOI222X1 U5408 (.IN1(sboxw[3]), .IN2(n6950), .IN3(n7090), .IN4(key[3]), .IN5(key[131])
          , .IN6(n6711), .QN(n3380));
   AOI222X1 U5409 (.IN1(n2924), .IN2(n7056), .IN3(n2921), .IN4(n7146), .IN5(n2923), .IN6(
          n7098), .QN(n3386));
   XOR2X1 U5410 (.IN1(n3387), .IN2(n7593), .Q(n2923));
   XOR2X1 U5411 (.IN1(n3387), .IN2(n7616), .Q(n2921));
   XOR3X1 U5412 (.IN1(prev_key0_reg[98]), .IN2(prev_key0_reg[66]), .IN3(n3388), .Q(n3387)
          );
   XNOR2X1 U5413 (.IN1(prev_key0_reg[2]), .IN2(prev_key0_reg[34]), .Q(n3388));
   XNOR3X1 U5414 (.IN1(prev_key1_reg[34]), .IN2(new_sboxw[26]), .IN3(n3389), .Q(n2924));
   XNOR3X1 U5415 (.IN1(sboxw[2]), .IN2(prev_key1_reg[98]), .IN3(prev_key1_reg[66]), .Q(
          n3389));
   AOI222X1 U5416 (.IN1(sboxw[2]), .IN2(n6950), .IN3(n7090), .IN4(key[2]), .IN5(key[130])
          , .IN6(n2945), .QN(n3385));
   AOI222X1 U5417 (.IN1(n2929), .IN2(n7056), .IN3(n2926), .IN4(n7146), .IN5(n2928), .IN6(
          n7098), .QN(n3391));
   XOR2X1 U5418 (.IN1(n3392), .IN2(n7592), .Q(n2928));
   XOR2X1 U5419 (.IN1(n3392), .IN2(n7615), .Q(n2926));
   XOR3X1 U5420 (.IN1(prev_key0_reg[97]), .IN2(prev_key0_reg[65]), .IN3(n3393), .Q(n3392)
          );
   XNOR2X1 U5421 (.IN1(prev_key0_reg[1]), .IN2(prev_key0_reg[33]), .Q(n3393));
   XNOR3X1 U5422 (.IN1(prev_key1_reg[33]), .IN2(new_sboxw[25]), .IN3(n3394), .Q(n2929));
   XNOR3X1 U5423 (.IN1(sboxw[1]), .IN2(prev_key1_reg[97]), .IN3(prev_key1_reg[65]), .Q(
          n3394));
   AOI222X1 U5424 (.IN1(sboxw[1]), .IN2(n6951), .IN3(n7090), .IN4(key[1]), .IN5(key[129])
          , .IN6(n6710), .QN(n3390));
   AO222X1 U5425 (.IN1(n6957), .IN2(key[255]), .IN3(prev_key1_reg[127]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[127]), .Q(n5473));
   AO222X1 U5426 (.IN1(n6958), .IN2(key[254]), .IN3(prev_key1_reg[126]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[126]), .Q(n5474));
   AO222X1 U5427 (.IN1(n6958), .IN2(key[253]), .IN3(prev_key1_reg[125]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[125]), .Q(n5475));
   AO222X1 U5428 (.IN1(n6960), .IN2(key[252]), .IN3(prev_key1_reg[124]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[124]), .Q(n5476));
   AO222X1 U5429 (.IN1(n6961), .IN2(key[251]), .IN3(prev_key1_reg[123]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[123]), .Q(n5477));
   AO222X1 U5430 (.IN1(n6959), .IN2(key[250]), .IN3(prev_key1_reg[122]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[122]), .Q(n5478));
   AO222X1 U5431 (.IN1(n6959), .IN2(key[249]), .IN3(prev_key1_reg[121]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[121]), .Q(n5479));
   AO222X1 U5432 (.IN1(n6960), .IN2(key[248]), .IN3(prev_key1_reg[120]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[120]), .Q(n5480));
   AO222X1 U5433 (.IN1(n6961), .IN2(key[247]), .IN3(prev_key1_reg[119]), .IN4(n6903), .IN5(
          n7023), .IN6(prev_key0_reg[119]), .Q(n5481));
   AO222X1 U5434 (.IN1(n6962), .IN2(key[246]), .IN3(prev_key1_reg[118]), .IN4(n6904), .IN5(
          n7023), .IN6(prev_key0_reg[118]), .Q(n5482));
   AO222X1 U5435 (.IN1(n6963), .IN2(key[245]), .IN3(prev_key1_reg[117]), .IN4(n6904), .IN5(
          n7023), .IN6(prev_key0_reg[117]), .Q(n5483));
   AO222X1 U5436 (.IN1(n6959), .IN2(key[244]), .IN3(prev_key1_reg[116]), .IN4(n6904), .IN5(
          n7023), .IN6(prev_key0_reg[116]), .Q(n5484));
   AO222X1 U5437 (.IN1(n6962), .IN2(key[243]), .IN3(prev_key1_reg[115]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[115]), .Q(n5485));
   AO222X1 U5438 (.IN1(n6963), .IN2(key[242]), .IN3(prev_key1_reg[114]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[114]), .Q(n5486));
   AO222X1 U5439 (.IN1(n6961), .IN2(key[241]), .IN3(prev_key1_reg[113]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[113]), .Q(n5487));
   AO222X1 U5440 (.IN1(n6962), .IN2(key[240]), .IN3(prev_key1_reg[112]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[112]), .Q(n5488));
   AO222X1 U5441 (.IN1(n6963), .IN2(key[239]), .IN3(prev_key1_reg[111]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[111]), .Q(n5489));
   AO222X1 U5442 (.IN1(n6964), .IN2(key[238]), .IN3(prev_key1_reg[110]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[110]), .Q(n5490));
   AO222X1 U5443 (.IN1(n6965), .IN2(key[237]), .IN3(prev_key1_reg[109]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[109]), .Q(n5491));
   AO222X1 U5444 (.IN1(n6957), .IN2(key[236]), .IN3(prev_key1_reg[108]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[108]), .Q(n5492));
   AO222X1 U5445 (.IN1(n6965), .IN2(key[235]), .IN3(prev_key1_reg[107]), .IN4(n6904), .IN5(
          n7024), .IN6(prev_key0_reg[107]), .Q(n5493));
   AO222X1 U5446 (.IN1(n6957), .IN2(key[234]), .IN3(prev_key1_reg[106]), .IN4(n6905), .IN5(
          n7024), .IN6(prev_key0_reg[106]), .Q(n5494));
   AO222X1 U5447 (.IN1(n6958), .IN2(key[233]), .IN3(prev_key1_reg[105]), .IN4(n6905), .IN5(
          n7024), .IN6(prev_key0_reg[105]), .Q(n5495));
   AO222X1 U5448 (.IN1(n6957), .IN2(key[232]), .IN3(prev_key1_reg[104]), .IN4(n6905), .IN5(
          n7024), .IN6(prev_key0_reg[104]), .Q(n5496));
   AO222X1 U5449 (.IN1(n6958), .IN2(key[231]), .IN3(prev_key1_reg[103]), .IN4(n6905), .IN5(
          n7025), .IN6(prev_key0_reg[103]), .Q(n5497));
   AO222X1 U5450 (.IN1(n6959), .IN2(key[230]), .IN3(prev_key1_reg[102]), .IN4(n6905), .IN5(
          n7025), .IN6(prev_key0_reg[102]), .Q(n5498));
   AO222X1 U5451 (.IN1(n6960), .IN2(key[229]), .IN3(prev_key1_reg[101]), .IN4(n6905), .IN5(
          n7025), .IN6(prev_key0_reg[101]), .Q(n5499));
   AO222X1 U5452 (.IN1(n6961), .IN2(key[228]), .IN3(prev_key1_reg[100]), .IN4(n6905), .IN5(
          n7025), .IN6(prev_key0_reg[100]), .Q(n5500));
   AO222X1 U5453 (.IN1(n6958), .IN2(key[227]), .IN3(prev_key1_reg[99]), .IN4(n6905), .IN5(
          n7025), .IN6(prev_key0_reg[99]), .Q(n5501));
   AO222X1 U5454 (.IN1(n6959), .IN2(key[226]), .IN3(prev_key1_reg[98]), .IN4(n6903), .IN5(
          n7025), .IN6(prev_key0_reg[98]), .Q(n5502));
   AO222X1 U5455 (.IN1(n6960), .IN2(key[225]), .IN3(prev_key1_reg[97]), .IN4(n6903), .IN5(
          n7025), .IN6(prev_key0_reg[97]), .Q(n5503));
   AO222X1 U5456 (.IN1(n6964), .IN2(key[224]), .IN3(prev_key1_reg[96]), .IN4(n6903), .IN5(
          n7025), .IN6(prev_key0_reg[96]), .Q(n5504));
   AO222X1 U5457 (.IN1(n6962), .IN2(key[223]), .IN3(prev_key1_reg[95]), .IN4(n6902), .IN5(
          n7025), .IN6(prev_key0_reg[95]), .Q(n5505));
   AO222X1 U5458 (.IN1(n6963), .IN2(key[222]), .IN3(prev_key1_reg[94]), .IN4(n6902), .IN5(
          n7025), .IN6(prev_key0_reg[94]), .Q(n5506));
   AO222X1 U5459 (.IN1(n6964), .IN2(key[221]), .IN3(prev_key1_reg[93]), .IN4(n6902), .IN5(
          n7025), .IN6(prev_key0_reg[93]), .Q(n5507));
   AO222X1 U5460 (.IN1(n6965), .IN2(key[220]), .IN3(prev_key1_reg[92]), .IN4(n6902), .IN5(
          n7025), .IN6(prev_key0_reg[92]), .Q(n5508));
   AO222X1 U5461 (.IN1(n6957), .IN2(key[219]), .IN3(prev_key1_reg[91]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[91]), .Q(n5509));
   AO222X1 U5462 (.IN1(n6964), .IN2(key[218]), .IN3(prev_key1_reg[90]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[90]), .Q(n5510));
   AO222X1 U5463 (.IN1(n6961), .IN2(key[217]), .IN3(prev_key1_reg[89]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[89]), .Q(n5511));
   AO222X1 U5464 (.IN1(n6962), .IN2(key[216]), .IN3(prev_key1_reg[88]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[88]), .Q(n5512));
   AO222X1 U5465 (.IN1(n6965), .IN2(key[215]), .IN3(prev_key1_reg[87]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[87]), .Q(n5513));
   AO222X1 U5466 (.IN1(n6958), .IN2(key[214]), .IN3(prev_key1_reg[86]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[86]), .Q(n5514));
   AO222X1 U5467 (.IN1(n6959), .IN2(key[213]), .IN3(prev_key1_reg[85]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[85]), .Q(n5515));
   AO222X1 U5468 (.IN1(n6960), .IN2(key[212]), .IN3(prev_key1_reg[84]), .IN4(n6902), .IN5(
          n7026), .IN6(prev_key0_reg[84]), .Q(n5516));
   AO222X1 U5469 (.IN1(n6961), .IN2(key[211]), .IN3(prev_key1_reg[83]), .IN4(n6901), .IN5(
          n7026), .IN6(prev_key0_reg[83]), .Q(n5517));
   AO222X1 U5470 (.IN1(n6962), .IN2(key[210]), .IN3(prev_key1_reg[82]), .IN4(n6901), .IN5(
          n7026), .IN6(prev_key0_reg[82]), .Q(n5518));
   AO222X1 U5471 (.IN1(n6965), .IN2(key[209]), .IN3(prev_key1_reg[81]), .IN4(n6901), .IN5(
          n7026), .IN6(prev_key0_reg[81]), .Q(n5519));
   AO222X1 U5472 (.IN1(n6963), .IN2(key[208]), .IN3(prev_key1_reg[80]), .IN4(n6901), .IN5(
          n7026), .IN6(prev_key0_reg[80]), .Q(n5520));
   AO222X1 U5473 (.IN1(n6964), .IN2(key[207]), .IN3(prev_key1_reg[79]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[79]), .Q(n5521));
   AO222X1 U5474 (.IN1(n6957), .IN2(key[206]), .IN3(prev_key1_reg[78]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[78]), .Q(n5522));
   AO222X1 U5475 (.IN1(n6963), .IN2(key[205]), .IN3(prev_key1_reg[77]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[77]), .Q(n5523));
   AO222X1 U5476 (.IN1(n6964), .IN2(key[204]), .IN3(prev_key1_reg[76]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[76]), .Q(n5524));
   AO222X1 U5477 (.IN1(n6965), .IN2(key[203]), .IN3(prev_key1_reg[75]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[75]), .Q(n5525));
   AO222X1 U5478 (.IN1(n6965), .IN2(key[202]), .IN3(prev_key1_reg[74]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[74]), .Q(n5526));
   AO222X1 U5479 (.IN1(n6957), .IN2(key[201]), .IN3(prev_key1_reg[73]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[73]), .Q(n5527));
   AO222X1 U5480 (.IN1(n6964), .IN2(key[200]), .IN3(prev_key1_reg[72]), .IN4(n6901), .IN5(
          n7027), .IN6(prev_key0_reg[72]), .Q(n5528));
   AO222X1 U5481 (.IN1(n6957), .IN2(key[199]), .IN3(prev_key1_reg[71]), .IN4(n6900), .IN5(
          n7027), .IN6(prev_key0_reg[71]), .Q(n5529));
   AO222X1 U5482 (.IN1(n6958), .IN2(key[198]), .IN3(prev_key1_reg[70]), .IN4(n6900), .IN5(
          n7027), .IN6(prev_key0_reg[70]), .Q(n5530));
   AO222X1 U5483 (.IN1(n6959), .IN2(key[197]), .IN3(prev_key1_reg[69]), .IN4(n6900), .IN5(
          n7027), .IN6(prev_key0_reg[69]), .Q(n5531));
   AO222X1 U5484 (.IN1(n6960), .IN2(key[196]), .IN3(prev_key1_reg[68]), .IN4(n6900), .IN5(
          n7027), .IN6(prev_key0_reg[68]), .Q(n5532));
   AO222X1 U5485 (.IN1(n6961), .IN2(key[195]), .IN3(prev_key1_reg[67]), .IN4(n6900), .IN5(
          n7028), .IN6(prev_key0_reg[67]), .Q(n5533));
   AO222X1 U5486 (.IN1(n6958), .IN2(key[194]), .IN3(prev_key1_reg[66]), .IN4(n6897), .IN5(
          n7028), .IN6(prev_key0_reg[66]), .Q(n5534));
   AO222X1 U5487 (.IN1(n6962), .IN2(key[193]), .IN3(prev_key1_reg[65]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[65]), .Q(n5535));
   AO222X1 U5488 (.IN1(n6963), .IN2(key[192]), .IN3(prev_key1_reg[64]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[64]), .Q(n5536));
   AO222X1 U5489 (.IN1(n6965), .IN2(key[191]), .IN3(prev_key1_reg[63]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[63]), .Q(n5537));
   AO222X1 U5490 (.IN1(n6962), .IN2(key[190]), .IN3(prev_key1_reg[62]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[62]), .Q(n5538));
   AO222X1 U5491 (.IN1(n6963), .IN2(key[189]), .IN3(prev_key1_reg[61]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[61]), .Q(n5539));
   AO222X1 U5492 (.IN1(n6964), .IN2(key[188]), .IN3(prev_key1_reg[60]), .IN4(n6900), .IN5(
          n7028), .IN6(prev_key0_reg[60]), .Q(n5540));
   AO222X1 U5493 (.IN1(n6965), .IN2(key[187]), .IN3(prev_key1_reg[59]), .IN4(n6899), .IN5(
          n7028), .IN6(prev_key0_reg[59]), .Q(n5541));
   AO222X1 U5494 (.IN1(n6957), .IN2(key[186]), .IN3(prev_key1_reg[58]), .IN4(n6897), .IN5(
          n7028), .IN6(prev_key0_reg[58]), .Q(n5542));
   AO222X1 U5495 (.IN1(n6959), .IN2(key[185]), .IN3(prev_key1_reg[57]), .IN4(n6897), .IN5(
          n7028), .IN6(prev_key0_reg[57]), .Q(n5543));
   AO222X1 U5496 (.IN1(n6964), .IN2(key[184]), .IN3(prev_key1_reg[56]), .IN4(n6900), .IN5(
          n7028), .IN6(prev_key0_reg[56]), .Q(n5544));
   AO222X1 U5497 (.IN1(n6965), .IN2(key[183]), .IN3(prev_key1_reg[55]), .IN4(n6899), .IN5(
          n7029), .IN6(prev_key0_reg[55]), .Q(n5545));
   AO222X1 U5498 (.IN1(n6957), .IN2(key[182]), .IN3(prev_key1_reg[54]), .IN4(n6897), .IN5(
          n7029), .IN6(prev_key0_reg[54]), .Q(n5546));
   AO222X1 U5499 (.IN1(n6958), .IN2(key[181]), .IN3(prev_key1_reg[53]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[53]), .Q(n5547));
   AO222X1 U5500 (.IN1(n6959), .IN2(key[180]), .IN3(prev_key1_reg[52]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[52]), .Q(n5548));
   AO222X1 U5501 (.IN1(n6960), .IN2(key[179]), .IN3(prev_key1_reg[51]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[51]), .Q(n5549));
   AO222X1 U5502 (.IN1(n6961), .IN2(key[178]), .IN3(prev_key1_reg[50]), .IN4(n6899), .IN5(
          n7029), .IN6(prev_key0_reg[50]), .Q(n5550));
   AO222X1 U5503 (.IN1(n6962), .IN2(key[177]), .IN3(prev_key1_reg[49]), .IN4(n6899), .IN5(
          n7029), .IN6(prev_key0_reg[49]), .Q(n5551));
   AO222X1 U5504 (.IN1(n6960), .IN2(key[176]), .IN3(prev_key1_reg[48]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[48]), .Q(n5552));
   AO222X1 U5505 (.IN1(n6957), .IN2(key[175]), .IN3(prev_key1_reg[47]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[47]), .Q(n5553));
   AO222X1 U5506 (.IN1(n6958), .IN2(key[174]), .IN3(prev_key1_reg[46]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[46]), .Q(n5554));
   AO222X1 U5507 (.IN1(n6958), .IN2(key[173]), .IN3(prev_key1_reg[45]), .IN4(n6898), .IN5(
          n7029), .IN6(prev_key0_reg[45]), .Q(n5555));
   AO222X1 U5508 (.IN1(n6963), .IN2(key[172]), .IN3(prev_key1_reg[44]), .IN4(n6899), .IN5(
          n7029), .IN6(prev_key0_reg[44]), .Q(n5556));
   AO222X1 U5509 (.IN1(n6964), .IN2(key[171]), .IN3(prev_key1_reg[43]), .IN4(n6900), .IN5(
          n7030), .IN6(prev_key0_reg[43]), .Q(n5557));
   AO222X1 U5510 (.IN1(n6965), .IN2(key[170]), .IN3(prev_key1_reg[42]), .IN4(n6899), .IN5(
          n7030), .IN6(prev_key0_reg[42]), .Q(n5558));
   AO222X1 U5511 (.IN1(n6957), .IN2(key[169]), .IN3(prev_key1_reg[41]), .IN4(n6898), .IN5(
          n7030), .IN6(prev_key0_reg[41]), .Q(n5559));
   AO222X1 U5512 (.IN1(n6958), .IN2(key[168]), .IN3(prev_key1_reg[40]), .IN4(n6898), .IN5(
          n7030), .IN6(prev_key0_reg[40]), .Q(n5560));
   AO222X1 U5513 (.IN1(n6961), .IN2(key[167]), .IN3(prev_key1_reg[39]), .IN4(n6900), .IN5(
          n7030), .IN6(prev_key0_reg[39]), .Q(n5561));
   AO222X1 U5514 (.IN1(n6959), .IN2(key[166]), .IN3(prev_key1_reg[38]), .IN4(n6898), .IN5(
          n7030), .IN6(prev_key0_reg[38]), .Q(n5562));
   AO222X1 U5515 (.IN1(n6960), .IN2(key[165]), .IN3(prev_key1_reg[37]), .IN4(n6898), .IN5(
          n7030), .IN6(prev_key0_reg[37]), .Q(n5563));
   AO222X1 U5516 (.IN1(n6959), .IN2(key[164]), .IN3(prev_key1_reg[36]), .IN4(n6898), .IN5(
          n7030), .IN6(prev_key0_reg[36]), .Q(n5564));
   AO222X1 U5517 (.IN1(n6959), .IN2(key[163]), .IN3(prev_key1_reg[35]), .IN4(n6899), .IN5(
          n7030), .IN6(prev_key0_reg[35]), .Q(n5565));
   AO222X1 U5518 (.IN1(n6960), .IN2(key[162]), .IN3(prev_key1_reg[34]), .IN4(n6895), .IN5(
          n7030), .IN6(prev_key0_reg[34]), .Q(n5566));
   AO222X1 U5519 (.IN1(n6961), .IN2(key[161]), .IN3(prev_key1_reg[33]), .IN4(n6896), .IN5(
          n7030), .IN6(prev_key0_reg[33]), .Q(n5567));
   AO222X1 U5520 (.IN1(n6962), .IN2(key[160]), .IN3(prev_key1_reg[32]), .IN4(n6896), .IN5(
          n7030), .IN6(prev_key0_reg[32]), .Q(n5568));
   AO222X1 U5521 (.IN1(n6963), .IN2(key[159]), .IN3(sboxw[31]), .IN4(n6896), .IN5(n7031), .
          IN6(prev_key0_reg[31]), .Q(n5569));
   AO222X1 U5522 (.IN1(n6961), .IN2(key[158]), .IN3(sboxw[30]), .IN4(n6896), .IN5(n7031), .
          IN6(prev_key0_reg[30]), .Q(n5570));
   AO222X1 U5523 (.IN1(n6965), .IN2(key[157]), .IN3(sboxw[29]), .IN4(n6896), .IN5(n7031), .
          IN6(prev_key0_reg[29]), .Q(n5571));
   AO222X1 U5524 (.IN1(n6957), .IN2(key[156]), .IN3(sboxw[28]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[28]), .Q(n5572));
   AO222X1 U5525 (.IN1(n6960), .IN2(key[155]), .IN3(sboxw[27]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[27]), .Q(n5573));
   AO222X1 U5526 (.IN1(n6964), .IN2(key[154]), .IN3(sboxw[26]), .IN4(n6897), .IN5(n7031), .
          IN6(prev_key0_reg[26]), .Q(n5574));
   AO222X1 U5527 (.IN1(n6965), .IN2(key[153]), .IN3(sboxw[25]), .IN4(n6896), .IN5(n7031), .
          IN6(prev_key0_reg[25]), .Q(n5575));
   AO222X1 U5528 (.IN1(n6957), .IN2(key[152]), .IN3(sboxw[24]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[24]), .Q(n5576));
   AO222X1 U5529 (.IN1(n6958), .IN2(key[151]), .IN3(sboxw[23]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[23]), .Q(n5577));
   AO222X1 U5530 (.IN1(n6959), .IN2(key[150]), .IN3(sboxw[22]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[22]), .Q(n5578));
   AO222X1 U5531 (.IN1(n6962), .IN2(key[149]), .IN3(sboxw[21]), .IN4(n6896), .IN5(n7031), .
          IN6(prev_key0_reg[21]), .Q(n5579));
   AO222X1 U5532 (.IN1(n6958), .IN2(key[148]), .IN3(sboxw[20]), .IN4(n6895), .IN5(n7031), .
          IN6(prev_key0_reg[20]), .Q(n5580));
   AO222X1 U5533 (.IN1(n6959), .IN2(key[147]), .IN3(sboxw[19]), .IN4(n6895), .IN5(n7032), .
          IN6(prev_key0_reg[19]), .Q(n5581));
   AO222X1 U5534 (.IN1(n6961), .IN2(key[146]), .IN3(sboxw[18]), .IN4(n6896), .IN5(n7032), .
          IN6(prev_key0_reg[18]), .Q(n5582));
   AO222X1 U5535 (.IN1(n6960), .IN2(key[145]), .IN3(sboxw[17]), .IN4(n6895), .IN5(n7032), .
          IN6(prev_key0_reg[17]), .Q(n5583));
   AO222X1 U5536 (.IN1(n6961), .IN2(key[144]), .IN3(sboxw[16]), .IN4(n6896), .IN5(n7032), .
          IN6(prev_key0_reg[16]), .Q(n5584));
   AO222X1 U5537 (.IN1(n6962), .IN2(key[143]), .IN3(sboxw[15]), .IN4(n6896), .IN5(n7032), .
          IN6(prev_key0_reg[15]), .Q(n5585));
   AO222X1 U5538 (.IN1(n6963), .IN2(key[142]), .IN3(sboxw[14]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[14]), .Q(n5586));
   AO222X1 U5539 (.IN1(n6964), .IN2(key[141]), .IN3(sboxw[13]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[13]), .Q(n5587));
   AO222X1 U5540 (.IN1(n6963), .IN2(key[140]), .IN3(sboxw[12]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[12]), .Q(n5588));
   AO222X1 U5541 (.IN1(n6960), .IN2(key[139]), .IN3(sboxw[11]), .IN4(n6895), .IN5(n7032), .
          IN6(prev_key0_reg[11]), .Q(n5589));
   AO222X1 U5542 (.IN1(n6961), .IN2(key[138]), .IN3(sboxw[10]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[10]), .Q(n5590));
   AO222X1 U5543 (.IN1(n6962), .IN2(key[137]), .IN3(sboxw[9]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[9]), .Q(n5591));
   AO222X1 U5544 (.IN1(n6965), .IN2(key[136]), .IN3(sboxw[8]), .IN4(n6897), .IN5(n7032), .
          IN6(prev_key0_reg[8]), .Q(n5592));
   AO222X1 U5545 (.IN1(n6957), .IN2(key[135]), .IN3(sboxw[7]), .IN4(n6895), .IN5(n7033), .
          IN6(prev_key0_reg[7]), .Q(n5593));
   AO222X1 U5546 (.IN1(n6958), .IN2(key[134]), .IN3(sboxw[6]), .IN4(n6895), .IN5(n7033), .
          IN6(prev_key0_reg[6]), .Q(n5594));
   AO222X1 U5547 (.IN1(n6959), .IN2(key[133]), .IN3(sboxw[5]), .IN4(n6896), .IN5(n7033), .
          IN6(prev_key0_reg[5]), .Q(n5595));
   AO222X1 U5548 (.IN1(n6960), .IN2(key[132]), .IN3(sboxw[4]), .IN4(n6896), .IN5(n7033), .
          IN6(prev_key0_reg[4]), .Q(n5596));
   AO222X1 U5549 (.IN1(n6964), .IN2(key[131]), .IN3(sboxw[3]), .IN4(n6897), .IN5(n7033), .
          IN6(prev_key0_reg[3]), .Q(n5597));
   AO222X1 U5550 (.IN1(n6962), .IN2(key[130]), .IN3(sboxw[2]), .IN4(n6900), .IN5(n7033), .
          IN6(prev_key0_reg[2]), .Q(n5598));
   AO222X1 U5551 (.IN1(n6963), .IN2(key[129]), .IN3(sboxw[1]), .IN4(n6900), .IN5(n7033), .
          IN6(prev_key0_reg[1]), .Q(n5599));
   AO222X1 U5552 (.IN1(n6963), .IN2(key[128]), .IN3(sboxw[0]), .IN4(n6900), .IN5(n7033), .
          IN6(prev_key0_reg[0]), .Q(n5600));
   AOI222X1 U5553 (.IN1(n2940), .IN2(n7056), .IN3(n2937), .IN4(n7146), .IN5(n2939), .IN6(
          n7098), .QN(n3399));
   XOR2X1 U5554 (.IN1(n3400), .IN2(n7591), .Q(n2939));
   XOR2X1 U5556 (.IN1(n3400), .IN2(n7614), .Q(n2937));
   XOR3X1 U5557 (.IN1(prev_key0_reg[96]), .IN2(prev_key0_reg[64]), .IN3(n3402), .Q(n3400)
          );
   XNOR2X1 U5558 (.IN1(prev_key0_reg[0]), .IN2(prev_key0_reg[32]), .Q(n3402));
   XNOR3X1 U5560 (.IN1(prev_key1_reg[32]), .IN2(new_sboxw[24]), .IN3(n3404), .Q(n2940));
   XNOR3X1 U5561 (.IN1(sboxw[0]), .IN2(prev_key1_reg[96]), .IN3(prev_key1_reg[64]), .Q(
          n3404));
   AOI222X1 U5562 (.IN1(sboxw[0]), .IN2(n6950), .IN3(n7090), .IN4(key[0]), .IN5(key[128])
          , .IN6(n6709), .QN(n3398));
   AO22X1 U5565 (.IN1(ready), .IN2(n3408), .IN3(key_mem_ctrl_reg[1]), .IN4(
          key_mem_ctrl_reg[0]), .Q(n5602));
   AO221X1 U5566 (.IN1(rcon_reg[6]), .IN2(n3410), .IN3(n3411), .IN4(rcon_reg[7]), .IN5(
          n3412), .Q(n5603));
   AO22X1 U5567 (.IN1(n3411), .IN2(rcon_reg[6]), .IN3(rcon_reg[5]), .IN4(n3410), .Q(n5604)
          );
   AO22X1 U5568 (.IN1(n3411), .IN2(rcon_reg[5]), .IN3(rcon_reg[4]), .IN4(n3410), .Q(n5605)
          );
   AO22X1 U5569 (.IN1(n3411), .IN2(rcon_reg[4]), .IN3(n3413), .IN4(n3410), .Q(n5606));
   XOR2X1 U5570 (.IN1(rcon_reg[7]), .IN2(rcon_reg[3]), .Q(n3413));
   AO221X1 U5571 (.IN1(n3414), .IN2(n3410), .IN3(n3411), .IN4(rcon_reg[3]), .IN5(n3412), .
          Q(n5607));
   XOR2X1 U5572 (.IN1(rcon_reg[7]), .IN2(rcon_reg[2]), .Q(n3414));
   AO221X1 U5573 (.IN1(rcon_reg[1]), .IN2(n3410), .IN3(n3411), .IN4(rcon_reg[2]), .IN5(
          n3412), .Q(n5608));
   AO221X1 U5574 (.IN1(rcon_reg[7]), .IN2(n3410), .IN3(n3411), .IN4(rcon_reg[0]), .IN5(
          n3412), .Q(n5609));
   AO22X1 U5575 (.IN1(n3411), .IN2(rcon_reg[1]), .IN3(n3415), .IN4(n3410), .Q(n5610));
   XOR2X1 U5576 (.IN1(rcon_reg[7]), .IN2(rcon_reg[0]), .Q(n3415));
   OR2X1 U5577 (.IN1(n3405), .IN2(n2933), .Q(n3410));
   NOR3X0 U5579 (.IN1(round_ctr_reg[2]), .IN2(round_ctr_reg[3]), .IN3(round_ctr_reg[1]), .
          QN(n3407));
   AO222X1 U5580 (.IN1(n2933), .IN2(n2935), .IN3(n2936), .IN4(n7581), .IN5(
          round_ctr_reg[3]), .IN6(n3416), .Q(n5611));
   AND3X1 U5581 (.IN1(round_ctr_reg[1]), .IN2(n2212), .IN3(round_ctr_reg[2]), .Q(n2935));
   AO22X1 U5582 (.IN1(round_ctr_reg[2]), .IN2(n3416), .IN3(n3417), .IN4(n2933), .Q(n5612)
          );
   AO21X1 U5583 (.IN1(n7581), .IN2(n2213), .IN3(n3418), .Q(n3416));
   AO22X1 U5584 (.IN1(round_ctr_reg[1]), .IN2(n3418), .IN3(n2933), .IN4(n2213), .Q(n5613)
          );
   AO21X1 U5585 (.IN1(n7581), .IN2(n2214), .IN3(n3419), .Q(n3418));
   AO22X1 U5586 (.IN1(n3419), .IN2(round_ctr_reg[0]), .IN3(n7581), .IN4(n2214), .Q(n5614)
          );
   AO221X1 U5590 (.IN1(n3423), .IN2(n7581), .IN3(key_mem_ctrl_reg[0]), .IN4(n2204), .IN5(
          n7582), .Q(n5616));
   AND4X1 U5594 (.IN1(n3425), .IN2(round_ctr_reg[3]), .IN3(round_ctr_reg[1]), .IN4(n2214)
          , .Q(n3423));
   SDFFARX1 \key_mem_reg[1][110]  (.D(n3682), .SI(n9548), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7469), .Q(\key_mem[1][110] ), .QN(n9547));
   SDFFARX1 \round_ctr_reg_reg[0]  (.D(n5614), .SI(n7625), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7495), .Q(round_ctr_reg[0]), .QN(n2214));
   SDFFARX1 \round_ctr_reg_reg[2]  (.D(n5612), .SI(n2213), .SE(test_se_buf_net7), .CLK(
          clk_buf_net7), .RSTB(n7495), .Q(round_ctr_reg[2]), .QN(n7624));
   SDFFARX1 \key_mem_ctrl_reg_reg[1]  (.D(n5615), .SI(key_mem_ctrl_reg[0]), .SE(
          test_se_buf_net7), .CLK(clk_buf_net7), .RSTB(n7495), .Q(key_mem_ctrl_reg[1]), .
          QN(n2242));
   NBUFFX4 U2191 (.INP(n6457), .Z(n6591));
   NBUFFX4 U2192 (.INP(n6450), .Z(n6502));
   NBUFFX4 U2197 (.INP(n6463), .Z(n6667));
   NBUFFX2 U2198 (.INP(n6462), .Z(n6651));
   NBUFFX2 U2199 (.INP(n6460), .Z(n6623));
   NBUFFX2 U2200 (.INP(n6455), .Z(n6563));
   NBUFFX2 U2201 (.INP(n6465), .Z(n6683));
   NBUFFX2 U2202 (.INP(n6452), .Z(n6518));
   NBUFFX2 U2203 (.INP(n6454), .Z(n6548));
   NBUFFX2 U2204 (.INP(n6460), .Z(n6622));
   NBUFFX2 U2205 (.INP(n6455), .Z(n6562));
   NBUFFX2 U2206 (.INP(n6465), .Z(n6682));
   NBUFFX2 U2207 (.INP(n6452), .Z(n6517));
   NBUFFX2 U2208 (.INP(n6458), .Z(n6608));
   NBUFFX2 U2209 (.INP(n6454), .Z(n6547));
   NBUFFX2 U2210 (.INP(n6461), .Z(n6638));
   NBUFFX2 U2211 (.INP(n6458), .Z(n6607));
   NBUFFX2 U2212 (.INP(n6453), .Z(n6533));
   NBUFFX2 U2213 (.INP(n6456), .Z(n6578));
   NBUFFX2 U2214 (.INP(n6455), .Z(n6561));
   NBUFFX2 U2215 (.INP(n6465), .Z(n6681));
   NBUFFX2 U2216 (.INP(n6452), .Z(n6516));
   NBUFFX2 U2217 (.INP(n6461), .Z(n6637));
   NBUFFX2 U2218 (.INP(n6453), .Z(n6532));
   NBUFFX2 U2219 (.INP(n6456), .Z(n6577));
   NBUFFX2 U2220 (.INP(n6454), .Z(n6546));
   NBUFFX2 U2221 (.INP(n6453), .Z(n6531));
   NBUFFX2 U2222 (.INP(n6456), .Z(n6576));
   NBUFFX2 U2223 (.INP(n6466), .Z(n6698));
   NBUFFX2 U2224 (.INP(n6466), .Z(n6697));
   NBUFFX2 U2225 (.INP(n6466), .Z(n6696));
   INVX0 U2226 (.INP(reset_n), .ZN(n7579));
   XNOR3X1 U2227 (.IN1(n3), .IN2(n1), .IN3(n2), .Q(n2654));
   XNOR2X1 U2228 (.IN1(prev_key1_reg[120]), .IN2(n7583), .Q(n2));
   NAND3X0 U2229 (.IN1(keylen), .IN2(n7581), .IN3(n3401), .QN(n3397));
   NBUFFX2 U2230 (.INP(n7556), .Z(n7313));
   NBUFFX2 U2231 (.INP(n7556), .Z(n7314));
   NBUFFX2 U2232 (.INP(n7556), .Z(n7315));
   NBUFFX2 U2233 (.INP(n7555), .Z(n7316));
   NBUFFX2 U2234 (.INP(n7555), .Z(n7317));
   NBUFFX2 U2235 (.INP(n7555), .Z(n7318));
   NBUFFX2 U2236 (.INP(n7554), .Z(n7319));
   NBUFFX2 U2237 (.INP(n7554), .Z(n7320));
   NBUFFX2 U2238 (.INP(n7554), .Z(n7321));
   NBUFFX2 U2239 (.INP(n7553), .Z(n7322));
   NBUFFX2 U2240 (.INP(n7553), .Z(n7323));
   NBUFFX2 U2241 (.INP(n7553), .Z(n7324));
   NBUFFX2 U2242 (.INP(n7552), .Z(n7325));
   NBUFFX2 U2243 (.INP(n7552), .Z(n7326));
   NBUFFX2 U2244 (.INP(n7552), .Z(n7327));
   NBUFFX2 U2245 (.INP(n7551), .Z(n7328));
   NBUFFX2 U2246 (.INP(n7551), .Z(n7329));
   NBUFFX2 U2247 (.INP(n7551), .Z(n7330));
   NBUFFX2 U2248 (.INP(n7550), .Z(n7331));
   NBUFFX2 U2249 (.INP(n7550), .Z(n7332));
   NBUFFX2 U2250 (.INP(n7550), .Z(n7333));
   NBUFFX2 U2251 (.INP(n7549), .Z(n7334));
   NBUFFX2 U2252 (.INP(n7549), .Z(n7335));
   NBUFFX2 U2253 (.INP(n7549), .Z(n7336));
   NBUFFX2 U2254 (.INP(n7548), .Z(n7337));
   NBUFFX2 U2255 (.INP(n7548), .Z(n7338));
   NBUFFX2 U2256 (.INP(n7548), .Z(n7339));
   NBUFFX2 U2257 (.INP(n7547), .Z(n7340));
   NBUFFX2 U2258 (.INP(n7547), .Z(n7341));
   NBUFFX2 U2259 (.INP(n7547), .Z(n7342));
   NBUFFX2 U2260 (.INP(n7546), .Z(n7343));
   NBUFFX2 U2261 (.INP(n7546), .Z(n7344));
   NBUFFX2 U2262 (.INP(n7546), .Z(n7345));
   NBUFFX2 U2263 (.INP(n7545), .Z(n7346));
   NBUFFX2 U2264 (.INP(n7545), .Z(n7347));
   NBUFFX2 U2265 (.INP(n7545), .Z(n7348));
   NBUFFX2 U2266 (.INP(n7544), .Z(n7349));
   NBUFFX2 U2267 (.INP(n7544), .Z(n7350));
   NBUFFX2 U2268 (.INP(n7544), .Z(n7351));
   NBUFFX2 U2269 (.INP(n7543), .Z(n7352));
   NBUFFX2 U2270 (.INP(n7543), .Z(n7353));
   NBUFFX2 U2271 (.INP(n7543), .Z(n7354));
   NBUFFX2 U2272 (.INP(n7542), .Z(n7355));
   NBUFFX2 U2273 (.INP(n7542), .Z(n7356));
   NBUFFX2 U2274 (.INP(n7542), .Z(n7357));
   NBUFFX2 U2275 (.INP(n7541), .Z(n7358));
   NBUFFX2 U2276 (.INP(n7541), .Z(n7359));
   NBUFFX2 U2277 (.INP(n7541), .Z(n7360));
   NBUFFX2 U2278 (.INP(n7540), .Z(n7361));
   NBUFFX2 U2279 (.INP(n7540), .Z(n7362));
   NBUFFX2 U2280 (.INP(n7540), .Z(n7363));
   NBUFFX2 U2281 (.INP(n7539), .Z(n7364));
   NBUFFX2 U2282 (.INP(n7539), .Z(n7365));
   NBUFFX2 U2283 (.INP(n7539), .Z(n7366));
   NBUFFX2 U2284 (.INP(n7538), .Z(n7367));
   NBUFFX2 U2285 (.INP(n7538), .Z(n7368));
   NBUFFX2 U2286 (.INP(n7538), .Z(n7369));
   NBUFFX2 U2287 (.INP(n7537), .Z(n7370));
   NBUFFX2 U2288 (.INP(n7537), .Z(n7371));
   NBUFFX2 U2289 (.INP(n7537), .Z(n7372));
   NBUFFX2 U2290 (.INP(n7536), .Z(n7373));
   NBUFFX2 U2291 (.INP(n7536), .Z(n7374));
   NBUFFX2 U2292 (.INP(n7536), .Z(n7375));
   NBUFFX2 U2293 (.INP(n7535), .Z(n7376));
   NBUFFX2 U2294 (.INP(n7535), .Z(n7377));
   NBUFFX2 U2295 (.INP(n7535), .Z(n7378));
   NBUFFX2 U2296 (.INP(n7534), .Z(n7379));
   NBUFFX2 U2297 (.INP(n7534), .Z(n7380));
   NBUFFX2 U2298 (.INP(n7534), .Z(n7381));
   NBUFFX2 U2299 (.INP(n7533), .Z(n7382));
   NBUFFX2 U2300 (.INP(n7533), .Z(n7383));
   NBUFFX2 U2301 (.INP(n7533), .Z(n7384));
   NBUFFX2 U2302 (.INP(n7532), .Z(n7385));
   NBUFFX2 U2303 (.INP(n7532), .Z(n7386));
   NBUFFX2 U2304 (.INP(n7532), .Z(n7387));
   NBUFFX2 U2305 (.INP(n7531), .Z(n7388));
   NBUFFX2 U2306 (.INP(n7531), .Z(n7389));
   NBUFFX2 U2307 (.INP(n7531), .Z(n7390));
   NBUFFX2 U2308 (.INP(n7530), .Z(n7391));
   NBUFFX2 U2309 (.INP(n7530), .Z(n7392));
   NBUFFX2 U2310 (.INP(n7530), .Z(n7393));
   NBUFFX2 U2311 (.INP(n7529), .Z(n7394));
   NBUFFX2 U2312 (.INP(n7529), .Z(n7395));
   NBUFFX2 U2313 (.INP(n7529), .Z(n7396));
   NBUFFX2 U2314 (.INP(n7528), .Z(n7397));
   NBUFFX2 U2315 (.INP(n7528), .Z(n7398));
   NBUFFX2 U2316 (.INP(n7528), .Z(n7399));
   NBUFFX2 U2317 (.INP(n7527), .Z(n7400));
   NBUFFX2 U2318 (.INP(n7527), .Z(n7401));
   NBUFFX2 U2319 (.INP(n7527), .Z(n7402));
   NBUFFX2 U2320 (.INP(n7526), .Z(n7403));
   NBUFFX2 U2321 (.INP(n7526), .Z(n7404));
   NBUFFX2 U2322 (.INP(n7526), .Z(n7405));
   NBUFFX2 U2323 (.INP(n7525), .Z(n7406));
   NBUFFX2 U2324 (.INP(n7525), .Z(n7407));
   NBUFFX2 U2325 (.INP(n7525), .Z(n7408));
   NBUFFX2 U2326 (.INP(n7524), .Z(n7409));
   NBUFFX2 U2327 (.INP(n7524), .Z(n7410));
   NBUFFX2 U2328 (.INP(n7524), .Z(n7411));
   NBUFFX2 U2329 (.INP(n7523), .Z(n7412));
   NBUFFX2 U2330 (.INP(n7523), .Z(n7413));
   NBUFFX2 U2331 (.INP(n7523), .Z(n7414));
   NBUFFX2 U2332 (.INP(n7522), .Z(n7415));
   NBUFFX2 U2333 (.INP(n7522), .Z(n7416));
   NBUFFX2 U2334 (.INP(n7522), .Z(n7417));
   NBUFFX2 U2335 (.INP(n7521), .Z(n7418));
   NBUFFX2 U2336 (.INP(n7521), .Z(n7419));
   NBUFFX2 U2337 (.INP(n7521), .Z(n7420));
   NBUFFX2 U2338 (.INP(n7520), .Z(n7421));
   NBUFFX2 U2339 (.INP(n7520), .Z(n7422));
   NBUFFX2 U2340 (.INP(n7520), .Z(n7423));
   NBUFFX2 U2341 (.INP(n7519), .Z(n7424));
   NBUFFX2 U2342 (.INP(n7519), .Z(n7425));
   NBUFFX2 U2343 (.INP(n7519), .Z(n7426));
   NBUFFX2 U2344 (.INP(n7518), .Z(n7427));
   NBUFFX2 U2345 (.INP(n7518), .Z(n7428));
   NBUFFX2 U2346 (.INP(n7518), .Z(n7429));
   NBUFFX2 U2347 (.INP(n7517), .Z(n7430));
   NBUFFX2 U2348 (.INP(n7517), .Z(n7431));
   NBUFFX2 U2349 (.INP(n7517), .Z(n7432));
   NBUFFX2 U2350 (.INP(n7516), .Z(n7433));
   NBUFFX2 U2351 (.INP(n7516), .Z(n7434));
   NBUFFX2 U2352 (.INP(n7516), .Z(n7435));
   NBUFFX2 U2353 (.INP(n7515), .Z(n7436));
   NBUFFX2 U2354 (.INP(n7515), .Z(n7437));
   NBUFFX2 U2355 (.INP(n7515), .Z(n7438));
   NBUFFX2 U2356 (.INP(n7514), .Z(n7439));
   NBUFFX2 U2357 (.INP(n7514), .Z(n7440));
   NBUFFX2 U2358 (.INP(n7514), .Z(n7441));
   NBUFFX2 U2359 (.INP(n7513), .Z(n7442));
   NBUFFX2 U2360 (.INP(n7513), .Z(n7443));
   NBUFFX2 U2361 (.INP(n7513), .Z(n7444));
   NBUFFX2 U2362 (.INP(n7512), .Z(n7445));
   NBUFFX2 U2363 (.INP(n7512), .Z(n7446));
   NBUFFX2 U2364 (.INP(n7512), .Z(n7447));
   NBUFFX2 U2365 (.INP(n7511), .Z(n7448));
   NBUFFX2 U2366 (.INP(n7511), .Z(n7449));
   NBUFFX2 U2367 (.INP(n7511), .Z(n7450));
   NBUFFX2 U2368 (.INP(n7510), .Z(n7451));
   NBUFFX2 U2369 (.INP(n7510), .Z(n7452));
   NBUFFX2 U2370 (.INP(n7510), .Z(n7453));
   NBUFFX2 U2371 (.INP(n7509), .Z(n7454));
   NBUFFX2 U2372 (.INP(n7509), .Z(n7455));
   NBUFFX2 U2373 (.INP(n7509), .Z(n7456));
   NBUFFX2 U2374 (.INP(n7508), .Z(n7457));
   NBUFFX2 U2375 (.INP(n7508), .Z(n7458));
   NBUFFX2 U2376 (.INP(n7508), .Z(n7459));
   NBUFFX2 U2377 (.INP(n7507), .Z(n7460));
   NBUFFX2 U2378 (.INP(n7507), .Z(n7461));
   NBUFFX2 U2379 (.INP(n7507), .Z(n7462));
   NBUFFX2 U2380 (.INP(n7506), .Z(n7463));
   NBUFFX2 U2381 (.INP(n7506), .Z(n7464));
   NBUFFX2 U2382 (.INP(n7506), .Z(n7465));
   NBUFFX2 U2383 (.INP(n7505), .Z(n7466));
   NBUFFX2 U2384 (.INP(n7505), .Z(n7467));
   NBUFFX2 U2385 (.INP(n7505), .Z(n7468));
   NBUFFX2 U2386 (.INP(n7504), .Z(n7470));
   NBUFFX2 U2387 (.INP(n7504), .Z(n7471));
   NBUFFX2 U2388 (.INP(n7503), .Z(n7472));
   NBUFFX2 U2389 (.INP(n7503), .Z(n7473));
   NBUFFX2 U2390 (.INP(n7503), .Z(n7474));
   NBUFFX2 U2391 (.INP(n7502), .Z(n7475));
   NBUFFX2 U2392 (.INP(n7502), .Z(n7476));
   NBUFFX2 U2393 (.INP(n7502), .Z(n7477));
   NBUFFX2 U2394 (.INP(n7501), .Z(n7478));
   NBUFFX2 U2395 (.INP(n7501), .Z(n7479));
   NBUFFX2 U2396 (.INP(n7501), .Z(n7480));
   NBUFFX2 U2397 (.INP(n7500), .Z(n7481));
   NBUFFX2 U2398 (.INP(n7500), .Z(n7482));
   NBUFFX2 U2399 (.INP(n7500), .Z(n7483));
   NBUFFX2 U2400 (.INP(n7499), .Z(n7484));
   NBUFFX2 U2401 (.INP(n7499), .Z(n7485));
   NBUFFX2 U2402 (.INP(n7499), .Z(n7486));
   NBUFFX2 U2403 (.INP(n7498), .Z(n7487));
   NBUFFX2 U2404 (.INP(n7498), .Z(n7488));
   NBUFFX2 U2405 (.INP(n7498), .Z(n7489));
   NBUFFX2 U2421 (.INP(n7497), .Z(n7490));
   NBUFFX2 U2455 (.INP(n7497), .Z(n7491));
   NBUFFX2 U2472 (.INP(n7497), .Z(n7492));
   NBUFFX2 U2560 (.INP(n7504), .Z(n7469));
   NBUFFX2 U2574 (.INP(n6941), .Z(n6930));
   NBUFFX2 U2642 (.INP(n6940), .Z(n6934));
   NBUFFX2 U2727 (.INP(n6940), .Z(n6935));
   NBUFFX2 U2761 (.INP(n6939), .Z(n6937));
   NBUFFX2 U2778 (.INP(n6941), .Z(n6931));
   NBUFFX2 U2795 (.INP(n6941), .Z(n6932));
   NBUFFX2 U2812 (.INP(n6940), .Z(n6933));
   NBUFFX2 U2931 (.INP(n6939), .Z(n6936));
   NBUFFX2 U2948 (.INP(n6939), .Z(n6938));
   NBUFFX2 U3543 (.INP(n6942), .Z(n6928));
   NBUFFX2 U3560 (.INP(n6942), .Z(n6929));
   NBUFFX2 U3594 (.INP(n7496), .Z(n7493));
   NBUFFX2 U3611 (.INP(n7496), .Z(n7494));
   NBUFFX2 U3628 (.INP(n7496), .Z(n7495));
   NBUFFX2 U3730 (.INP(n7557), .Z(n7556));
   NBUFFX2 U3866 (.INP(n7557), .Z(n7555));
   NBUFFX2 U3883 (.INP(n7557), .Z(n7554));
   NBUFFX2 U3934 (.INP(n7558), .Z(n7553));
   NBUFFX2 U4019 (.INP(n7558), .Z(n7552));
   NBUFFX2 U4274 (.INP(n7558), .Z(n7551));
   NBUFFX2 U4359 (.INP(n7559), .Z(n7550));
   NBUFFX2 U4410 (.INP(n7559), .Z(n7549));
   NBUFFX2 U4427 (.INP(n7559), .Z(n7548));
   NBUFFX2 U4478 (.INP(n7560), .Z(n7547));
   NBUFFX2 U4512 (.INP(n7560), .Z(n7546));
   NBUFFX2 U4563 (.INP(n7560), .Z(n7545));
   NBUFFX2 U4571 (.INP(n7561), .Z(n7544));
   NBUFFX2 U4573 (.INP(n7561), .Z(n7543));
   NBUFFX2 U4577 (.INP(n7561), .Z(n7542));
   NBUFFX2 U4579 (.INP(n7562), .Z(n7541));
   NBUFFX2 U4581 (.INP(n7562), .Z(n7540));
   NBUFFX2 U4583 (.INP(n7562), .Z(n7539));
   NBUFFX2 U4585 (.INP(n7563), .Z(n7538));
   NBUFFX2 U4587 (.INP(n7563), .Z(n7537));
   NBUFFX2 U4588 (.INP(n7563), .Z(n7536));
   NBUFFX2 U4592 (.INP(n7564), .Z(n7535));
   NBUFFX2 U4640 (.INP(n7564), .Z(n7534));
   NBUFFX2 U4809 (.INP(n7564), .Z(n7533));
   NBUFFX2 U4850 (.INP(n7565), .Z(n7532));
   NBUFFX2 U4853 (.INP(n7565), .Z(n7531));
   NBUFFX2 U4862 (.INP(n7565), .Z(n7530));
   NBUFFX2 U4865 (.INP(n7566), .Z(n7529));
   NBUFFX2 U4880 (.INP(n7566), .Z(n7528));
   NBUFFX2 U4883 (.INP(n7566), .Z(n7527));
   NBUFFX2 U4886 (.INP(n7567), .Z(n7526));
   NBUFFX2 U4889 (.INP(n7567), .Z(n7525));
   NBUFFX2 U4899 (.INP(n7567), .Z(n7524));
   NBUFFX2 U4911 (.INP(n7568), .Z(n7523));
   NBUFFX2 U4929 (.INP(n7568), .Z(n7522));
   NBUFFX2 U4935 (.INP(n7568), .Z(n7521));
   NBUFFX2 U4998 (.INP(n7569), .Z(n7520));
   NBUFFX2 U4999 (.INP(n7569), .Z(n7519));
   NBUFFX2 U5075 (.INP(n7569), .Z(n7518));
   NBUFFX2 U5076 (.INP(n7570), .Z(n7517));
   NBUFFX2 U5237 (.INP(n7570), .Z(n7516));
   NBUFFX2 U5238 (.INP(n7570), .Z(n7515));
   NBUFFX2 U5310 (.INP(n7571), .Z(n7514));
   NBUFFX2 U5311 (.INP(n7571), .Z(n7513));
   NBUFFX2 U5326 (.INP(n7571), .Z(n7512));
   NBUFFX2 U5327 (.INP(n7572), .Z(n7511));
   NBUFFX2 U5350 (.INP(n7572), .Z(n7510));
   NBUFFX2 U5351 (.INP(n7572), .Z(n7509));
   NBUFFX2 U5555 (.INP(n7573), .Z(n7508));
   NBUFFX2 U5559 (.INP(n7573), .Z(n7507));
   NBUFFX2 U5563 (.INP(n7573), .Z(n7506));
   NBUFFX2 U5564 (.INP(n7574), .Z(n7505));
   NBUFFX2 U5578 (.INP(n7574), .Z(n7504));
   NBUFFX2 U5587 (.INP(n7574), .Z(n7503));
   NBUFFX2 U5588 (.INP(n7575), .Z(n7502));
   NBUFFX2 U5589 (.INP(n7575), .Z(n7501));
   NBUFFX2 U5591 (.INP(n7575), .Z(n7500));
   NBUFFX2 U5592 (.INP(n7576), .Z(n7499));
   NBUFFX2 U5593 (.INP(n7576), .Z(n7498));
   NBUFFX2 U5595 (.INP(n7576), .Z(n7497));
   NBUFFX2 U5596 (.INP(n6593), .Z(n6589));
   NBUFFX2 U5597 (.INP(n6488), .Z(n6484));
   NBUFFX2 U5598 (.INP(n6592), .Z(n6586));
   NBUFFX2 U5599 (.INP(n6487), .Z(n6481));
   NBUFFX2 U5600 (.INP(n6503), .Z(n6499));
   NBUFFX2 U5601 (.INP(n6668), .Z(n6664));
   NBUFFX2 U5602 (.INP(n6593), .Z(n6588));
   NBUFFX2 U5603 (.INP(n6488), .Z(n6483));
   NBUFFX2 U5604 (.INP(n6502), .Z(n6496));
   NBUFFX2 U5605 (.INP(n6667), .Z(n6661));
   NBUFFX2 U5606 (.INP(n6503), .Z(n6498));
   NBUFFX2 U5607 (.INP(n6668), .Z(n6663));
   NBUFFX2 U5608 (.INP(n6591), .Z(n6583));
   NBUFFX2 U5609 (.INP(n6486), .Z(n6478));
   NBUFFX2 U5610 (.INP(n6623), .Z(n6619));
   NBUFFX2 U5611 (.INP(n6591), .Z(n6582));
   NBUFFX2 U5612 (.INP(n6563), .Z(n6559));
   NBUFFX2 U5613 (.INP(n6683), .Z(n6679));
   NBUFFX2 U5614 (.INP(n6486), .Z(n6477));
   NBUFFX2 U5615 (.INP(n6518), .Z(n6514));
   NBUFFX2 U5616 (.INP(n6592), .Z(n6584));
   NBUFFX2 U5617 (.INP(n6487), .Z(n6479));
   NBUFFX2 U5618 (.INP(n6622), .Z(n6616));
   NBUFFX2 U5619 (.INP(n6548), .Z(n6544));
   NBUFFX2 U5620 (.INP(n6562), .Z(n6556));
   NBUFFX2 U5621 (.INP(n6682), .Z(n6676));
   NBUFFX2 U5622 (.INP(n6517), .Z(n6511));
   NBUFFX2 U5623 (.INP(n6501), .Z(n6493));
   NBUFFX2 U5624 (.INP(n6666), .Z(n6658));
   NBUFFX2 U5625 (.INP(n6501), .Z(n6492));
   NBUFFX2 U5626 (.INP(n6666), .Z(n6657));
   NBUFFX2 U5627 (.INP(n6502), .Z(n6494));
   NBUFFX2 U5628 (.INP(n6623), .Z(n6618));
   NBUFFX2 U5629 (.INP(n6667), .Z(n6659));
   NBUFFX2 U5630 (.INP(n6563), .Z(n6558));
   NBUFFX2 U5631 (.INP(n6547), .Z(n6541));
   NBUFFX2 U5632 (.INP(n6683), .Z(n6678));
   NBUFFX2 U5633 (.INP(n6518), .Z(n6513));
   NBUFFX2 U5634 (.INP(n6651), .Z(n6643));
   NBUFFX2 U5635 (.INP(n6638), .Z(n6634));
   NBUFFX2 U5636 (.INP(n6548), .Z(n6543));
   NBUFFX2 U5637 (.INP(n6533), .Z(n6529));
   NBUFFX2 U5638 (.INP(n6578), .Z(n6574));
   NBUFFX2 U5639 (.INP(n6651), .Z(n6642));
   NBUFFX2 U5640 (.INP(n6637), .Z(n6631));
   NBUFFX2 U5641 (.INP(n6532), .Z(n6526));
   NBUFFX2 U5642 (.INP(n6577), .Z(n6571));
   NBUFFX2 U5643 (.INP(n6638), .Z(n6633));
   NBUFFX2 U5644 (.INP(n6533), .Z(n6528));
   NBUFFX2 U5645 (.INP(n6578), .Z(n6573));
   NBUFFX2 U5646 (.INP(n6621), .Z(n6613));
   NBUFFX2 U5647 (.INP(n6591), .Z(n6581));
   NBUFFX2 U5648 (.INP(n6592), .Z(n6585));
   NBUFFX2 U5649 (.INP(n6561), .Z(n6553));
   NBUFFX2 U5650 (.INP(n6681), .Z(n6673));
   NBUFFX2 U5651 (.INP(n6486), .Z(n6476));
   NBUFFX2 U5652 (.INP(n6516), .Z(n6508));
   NBUFFX2 U5653 (.INP(n6487), .Z(n6480));
   NBUFFX2 U5654 (.INP(n6621), .Z(n6612));
   NBUFFX2 U5655 (.INP(n6561), .Z(n6552));
   NBUFFX2 U5656 (.INP(n6681), .Z(n6672));
   NBUFFX2 U5657 (.INP(n6516), .Z(n6507));
   NBUFFX2 U5658 (.INP(n6622), .Z(n6614));
   NBUFFX2 U5659 (.INP(n6562), .Z(n6554));
   NBUFFX2 U5660 (.INP(n6682), .Z(n6674));
   NBUFFX2 U5661 (.INP(n6517), .Z(n6509));
   NBUFFX2 U5662 (.INP(n6546), .Z(n6538));
   NBUFFX2 U5663 (.INP(n6593), .Z(n6587));
   NBUFFX2 U5664 (.INP(n6546), .Z(n6537));
   NBUFFX2 U5665 (.INP(n6488), .Z(n6482));
   NBUFFX2 U5666 (.INP(n6501), .Z(n6491));
   NBUFFX2 U5667 (.INP(n6502), .Z(n6495));
   NBUFFX2 U5668 (.INP(n6547), .Z(n6539));
   NBUFFX2 U5669 (.INP(n6666), .Z(n6656));
   NBUFFX2 U5670 (.INP(n6667), .Z(n6660));
   NBUFFX2 U5671 (.INP(n6608), .Z(n6604));
   NBUFFX2 U5672 (.INP(n6636), .Z(n6628));
   NBUFFX2 U5673 (.INP(n6503), .Z(n6497));
   NBUFFX2 U5674 (.INP(n6531), .Z(n6523));
   NBUFFX2 U5675 (.INP(n6576), .Z(n6568));
   NBUFFX2 U5676 (.INP(n6668), .Z(n6662));
   NBUFFX2 U5677 (.INP(n6607), .Z(n6601));
   NBUFFX2 U5678 (.INP(n6651), .Z(n6641));
   NBUFFX2 U5679 (.INP(n6636), .Z(n6627));
   NBUFFX2 U5680 (.INP(n6531), .Z(n6522));
   NBUFFX2 U5681 (.INP(n6576), .Z(n6567));
   NBUFFX2 U5682 (.INP(n6637), .Z(n6629));
   NBUFFX2 U5683 (.INP(n6532), .Z(n6524));
   NBUFFX2 U5684 (.INP(n6577), .Z(n6569));
   NBUFFX2 U5685 (.INP(n6608), .Z(n6603));
   NBUFFX2 U5686 (.INP(n6590), .Z(n6580));
   NBUFFX2 U5687 (.INP(n6485), .Z(n6475));
   NBUFFX2 U5688 (.INP(n6621), .Z(n6611));
   NBUFFX2 U5689 (.INP(n6622), .Z(n6615));
   NBUFFX2 U5690 (.INP(n6561), .Z(n6551));
   NBUFFX2 U5691 (.INP(n6681), .Z(n6671));
   NBUFFX2 U5692 (.INP(n6562), .Z(n6555));
   NBUFFX2 U5693 (.INP(n6682), .Z(n6675));
   NBUFFX2 U5694 (.INP(n6516), .Z(n6506));
   NBUFFX2 U5695 (.INP(n6517), .Z(n6510));
   NBUFFX2 U5696 (.INP(n6500), .Z(n6490));
   NBUFFX2 U5697 (.INP(n6665), .Z(n6655));
   NBUFFX2 U5698 (.INP(n6546), .Z(n6536));
   NBUFFX2 U5699 (.INP(n6547), .Z(n6540));
   NBUFFX2 U5700 (.INP(n6623), .Z(n6617));
   NBUFFX2 U5701 (.INP(n6563), .Z(n6557));
   NBUFFX2 U5702 (.INP(n6590), .Z(n6579));
   NBUFFX2 U5703 (.INP(n6683), .Z(n6677));
   NBUFFX2 U5704 (.INP(n6518), .Z(n6512));
   NBUFFX2 U5705 (.INP(n6485), .Z(n6474));
   NBUFFX2 U5706 (.INP(n6606), .Z(n6598));
   NBUFFX2 U5707 (.INP(n6650), .Z(n6640));
   NBUFFX2 U5708 (.INP(n6606), .Z(n6597));
   NBUFFX2 U5709 (.INP(n6548), .Z(n6542));
   NBUFFX2 U5710 (.INP(n6500), .Z(n6489));
   NBUFFX2 U5711 (.INP(n6607), .Z(n6599));
   NBUFFX2 U5712 (.INP(n6698), .Z(n6694));
   NBUFFX2 U5713 (.INP(n6665), .Z(n6654));
   NBUFFX2 U5714 (.INP(n6636), .Z(n6626));
   NBUFFX2 U5715 (.INP(n6637), .Z(n6630));
   NBUFFX2 U5716 (.INP(n6531), .Z(n6521));
   NBUFFX2 U5717 (.INP(n6576), .Z(n6566));
   NBUFFX2 U5718 (.INP(n6532), .Z(n6525));
   NBUFFX2 U5719 (.INP(n6577), .Z(n6570));
   NBUFFX2 U5720 (.INP(n6697), .Z(n6691));
   NBUFFX2 U5721 (.INP(n6638), .Z(n6632));
   NBUFFX2 U5722 (.INP(n6620), .Z(n6610));
   NBUFFX2 U5723 (.INP(n6533), .Z(n6527));
   NBUFFX2 U5724 (.INP(n6578), .Z(n6572));
   NBUFFX2 U5725 (.INP(n6560), .Z(n6550));
   NBUFFX2 U5726 (.INP(n6680), .Z(n6670));
   NBUFFX2 U5727 (.INP(n6698), .Z(n6693));
   NBUFFX2 U5728 (.INP(n6515), .Z(n6505));
   NBUFFX2 U5729 (.INP(n6650), .Z(n6639));
   NBUFFX2 U5730 (.INP(n6545), .Z(n6535));
   NBUFFX2 U5731 (.INP(n6635), .Z(n6625));
   NBUFFX2 U5732 (.INP(n6530), .Z(n6520));
   NBUFFX2 U5733 (.INP(n6575), .Z(n6565));
   NBUFFX2 U5734 (.INP(n6606), .Z(n6596));
   NBUFFX2 U5735 (.INP(n6620), .Z(n6609));
   NBUFFX2 U5736 (.INP(n6607), .Z(n6600));
   NBUFFX2 U5737 (.INP(n6560), .Z(n6549));
   NBUFFX2 U5738 (.INP(n6680), .Z(n6669));
   NBUFFX2 U5739 (.INP(n6515), .Z(n6504));
   NBUFFX2 U5740 (.INP(n6696), .Z(n6688));
   NBUFFX2 U5741 (.INP(n6696), .Z(n6687));
   NBUFFX2 U5742 (.INP(n6697), .Z(n6689));
   NBUFFX2 U5743 (.INP(n6545), .Z(n6534));
   NBUFFX2 U5744 (.INP(n6608), .Z(n6602));
   NBUFFX2 U5745 (.INP(n6635), .Z(n6624));
   NBUFFX2 U5746 (.INP(n6575), .Z(n6564));
   NBUFFX2 U5747 (.INP(n6530), .Z(n6519));
   NBUFFX2 U5748 (.INP(n6605), .Z(n6595));
   NBUFFX2 U5749 (.INP(n6696), .Z(n6686));
   NBUFFX2 U5750 (.INP(n6697), .Z(n6690));
   NBUFFX2 U5751 (.INP(n6605), .Z(n6594));
   NBUFFX2 U5752 (.INP(n6698), .Z(n6692));
   NBUFFX2 U5753 (.INP(n6695), .Z(n6685));
   NBUFFX2 U5754 (.INP(n6695), .Z(n6684));
   DELLN1X2 U5755 (.INP(n6653), .Z(n6649));
   DELLN1X2 U5756 (.INP(n6652), .Z(n6646));
   DELLN1X2 U5757 (.INP(n6653), .Z(n6648));
   DELLN1X2 U5758 (.INP(n6652), .Z(n6644));
   DELLN1X2 U5759 (.INP(n6652), .Z(n6645));
   DELLN1X2 U5760 (.INP(n6653), .Z(n6647));
   NBUFFX2 U5761 (.INP(n7035), .Z(n7030));
   NBUFFX2 U5762 (.INP(n7035), .Z(n7028));
   NBUFFX2 U5763 (.INP(n7036), .Z(n7027));
   NBUFFX2 U5764 (.INP(n7036), .Z(n7026));
   NBUFFX2 U5765 (.INP(n7036), .Z(n7025));
   NBUFFX2 U5766 (.INP(n7035), .Z(n7029));
   NBUFFX2 U5767 (.INP(n7037), .Z(n7024));
   NBUFFX2 U5768 (.INP(n7037), .Z(n7023));
   NBUFFX2 U5769 (.INP(n7310), .Z(n6941));
   NBUFFX2 U5770 (.INP(n7310), .Z(n6940));
   NBUFFX2 U5771 (.INP(n7310), .Z(n6939));
   NBUFFX2 U5772 (.INP(n6891), .Z(n6896));
   NBUFFX2 U5773 (.INP(n6892), .Z(n6899));
   NBUFFX2 U5774 (.INP(n6891), .Z(n6897));
   NBUFFX2 U5775 (.INP(n6892), .Z(n6900));
   NBUFFX2 U5776 (.INP(n6893), .Z(n6901));
   NBUFFX2 U5777 (.INP(n6893), .Z(n6902));
   NBUFFX2 U5778 (.INP(n6893), .Z(n6903));
   NBUFFX2 U5779 (.INP(n6891), .Z(n6895));
   NBUFFX2 U5780 (.INP(n6892), .Z(n6898));
   NBUFFX2 U5781 (.INP(n7310), .Z(n6942));
   NBUFFX2 U5782 (.INP(n6894), .Z(n6904));
   NBUFFX2 U5783 (.INP(n6894), .Z(n6905));
   NBUFFX2 U5784 (.INP(n7034), .Z(n7032));
   NBUFFX2 U5785 (.INP(n7034), .Z(n7031));
   NBUFFX2 U5786 (.INP(n7034), .Z(n7033));
   NBUFFX2 U5787 (.INP(n7577), .Z(n7557));
   NBUFFX2 U5788 (.INP(n7577), .Z(n7558));
   NBUFFX2 U5789 (.INP(n7566), .Z(n7559));
   NBUFFX2 U5790 (.INP(n7529), .Z(n7560));
   NBUFFX2 U5791 (.INP(n7528), .Z(n7561));
   NBUFFX2 U5792 (.INP(n7527), .Z(n7562));
   NBUFFX2 U5793 (.INP(n7567), .Z(n7563));
   NBUFFX2 U5794 (.INP(n7526), .Z(n7564));
   NBUFFX2 U5795 (.INP(n7525), .Z(n7565));
   NBUFFX2 U5796 (.INP(n7578), .Z(n7566));
   NBUFFX2 U5797 (.INP(n7578), .Z(n7567));
   NBUFFX2 U5798 (.INP(n7578), .Z(n7568));
   NBUFFX2 U5799 (.INP(n7578), .Z(n7569));
   NBUFFX2 U5800 (.INP(n7578), .Z(n7570));
   NBUFFX2 U5801 (.INP(n7578), .Z(n7571));
   NBUFFX2 U5802 (.INP(n7578), .Z(n7572));
   NBUFFX2 U5803 (.INP(n7578), .Z(n7573));
   NBUFFX2 U5804 (.INP(n7578), .Z(n7574));
   NBUFFX2 U5805 (.INP(n7578), .Z(n7575));
   NBUFFX2 U5806 (.INP(n7578), .Z(n7576));
   NBUFFX2 U5807 (.INP(n7577), .Z(n7496));
   NBUFFX2 U5808 (.INP(n7578), .Z(n7577));
   DELLN1X2 U5809 (.INP(n6457), .Z(n6593));
   DELLN1X2 U5810 (.INP(n6449), .Z(n6488));
   DELLN1X2 U5811 (.INP(n6457), .Z(n6592));
   DELLN1X2 U5812 (.INP(n6449), .Z(n6487));
   DELLN1X2 U5813 (.INP(n6450), .Z(n6503));
   DELLN1X2 U5814 (.INP(n6463), .Z(n6668));
   NBUFFX2 U5815 (.INP(n6449), .Z(n6486));
   NBUFFX2 U5816 (.INP(n6450), .Z(n6501));
   NBUFFX2 U5817 (.INP(n6463), .Z(n6666));
   NBUFFX2 U5818 (.INP(n6460), .Z(n6621));
   NBUFFX2 U5819 (.INP(n6461), .Z(n6636));
   NBUFFX2 U5820 (.INP(n6457), .Z(n6590));
   NBUFFX2 U5821 (.INP(n6449), .Z(n6485));
   NBUFFX2 U5822 (.INP(n6450), .Z(n6500));
   NBUFFX2 U5823 (.INP(n6463), .Z(n6665));
   NBUFFX2 U5824 (.INP(n6458), .Z(n6606));
   NBUFFX2 U5825 (.INP(n6462), .Z(n6650));
   NBUFFX2 U5826 (.INP(n6460), .Z(n6620));
   NBUFFX2 U5827 (.INP(n6455), .Z(n6560));
   NBUFFX2 U5828 (.INP(n6465), .Z(n6680));
   NBUFFX2 U5829 (.INP(n6452), .Z(n6515));
   NBUFFX2 U5830 (.INP(n6454), .Z(n6545));
   NBUFFX2 U5831 (.INP(n6461), .Z(n6635));
   NBUFFX2 U5832 (.INP(n6456), .Z(n6575));
   NBUFFX2 U5833 (.INP(n6453), .Z(n6530));
   NBUFFX2 U5834 (.INP(n6458), .Z(n6605));
   NBUFFX2 U5835 (.INP(n6466), .Z(n6695));
   NBUFFX2 U5836 (.INP(n7069), .Z(n7087));
   NBUFFX2 U5837 (.INP(n7069), .Z(n7086));
   NBUFFX2 U5838 (.INP(n7068), .Z(n7085));
   NBUFFX2 U5839 (.INP(n7068), .Z(n7084));
   NBUFFX2 U5840 (.INP(n7068), .Z(n7083));
   NBUFFX2 U5841 (.INP(n7069), .Z(n7088));
   NBUFFX2 U5842 (.INP(n3396), .Z(n7035));
   NBUFFX2 U5843 (.INP(n3396), .Z(n7036));
   NBUFFX2 U5844 (.INP(n7070), .Z(n7089));
   NBUFFX2 U5845 (.INP(n7610), .Z(n6700));
   NBUFFX2 U5846 (.INP(n7610), .Z(n6699));
   NBUFFX2 U5847 (.INP(n7610), .Z(n6701));
   NBUFFX2 U5848 (.INP(n7070), .Z(n7090));
   NBUFFX2 U5849 (.INP(n7059), .Z(n7048));
   NBUFFX2 U5850 (.INP(n3396), .Z(n7037));
   NBUFFX2 U5851 (.INP(n7060), .Z(n7047));
   NBUFFX2 U5852 (.INP(n7060), .Z(n7046));
   NBUFFX2 U5853 (.INP(n7060), .Z(n7045));
   NBUFFX2 U5854 (.INP(n7061), .Z(n7044));
   NBUFFX2 U5855 (.INP(n7061), .Z(n7043));
   NBUFFX2 U5856 (.INP(n7061), .Z(n7042));
   NBUFFX2 U5857 (.INP(n7062), .Z(n7041));
   NBUFFX2 U5858 (.INP(n7062), .Z(n7040));
   NBUFFX2 U5859 (.INP(n7062), .Z(n7039));
   NBUFFX2 U5860 (.INP(n7057), .Z(n7055));
   NBUFFX2 U5861 (.INP(n7057), .Z(n7054));
   NBUFFX2 U5862 (.INP(n7058), .Z(n7053));
   NBUFFX2 U5863 (.INP(n7058), .Z(n7052));
   NBUFFX2 U5864 (.INP(n7058), .Z(n7051));
   NBUFFX2 U5865 (.INP(n7059), .Z(n7050));
   NBUFFX2 U5866 (.INP(n7059), .Z(n7049));
   NBUFFX2 U5867 (.INP(n7580), .Z(n6891));
   NBUFFX2 U5868 (.INP(n7580), .Z(n6892));
   NBUFFX2 U5869 (.INP(n7580), .Z(n6893));
   NBUFFX2 U5870 (.INP(n7057), .Z(n7056));
   NBUFFX2 U5871 (.INP(n7580), .Z(n6894));
   NBUFFX2 U5872 (.INP(n2944), .Z(n6944));
   NBUFFX2 U5873 (.INP(n7067), .Z(n7081));
   NBUFFX2 U5874 (.INP(n7067), .Z(n7080));
   NBUFFX2 U5875 (.INP(n7066), .Z(n7079));
   NBUFFX2 U5876 (.INP(n7065), .Z(n7075));
   NBUFFX2 U5877 (.INP(n7064), .Z(n7072));
   NBUFFX2 U5878 (.INP(n7064), .Z(n7071));
   NBUFFX2 U5879 (.INP(n7066), .Z(n7078));
   NBUFFX2 U5880 (.INP(n7066), .Z(n7077));
   NBUFFX2 U5881 (.INP(n7065), .Z(n7076));
   NBUFFX2 U5882 (.INP(n7065), .Z(n7074));
   NBUFFX2 U5883 (.INP(n7064), .Z(n7073));
   NBUFFX2 U5884 (.INP(n7067), .Z(n7082));
   NBUFFX2 U5885 (.INP(n2944), .Z(n6946));
   NBUFFX2 U5886 (.INP(n2944), .Z(n6945));
   NBUFFX2 U5887 (.INP(n2944), .Z(n6948));
   NBUFFX2 U5888 (.INP(n2944), .Z(n6947));
   NBUFFX2 U5889 (.INP(n2944), .Z(n6949));
   NBUFFX2 U5890 (.INP(n3396), .Z(n7034));
   INVX0 U5891 (.INP(n7579), .ZN(n7578));
   NBUFFX2 U5892 (.INP(n7122), .Z(n7136));
   NBUFFX2 U5893 (.INP(n2297), .Z(n7069));
   NBUFFX2 U5894 (.INP(n2297), .Z(n7068));
   INVX0 U5895 (.INP(new_sboxw[22]), .ZN(n7605));
   NBUFFX2 U5896 (.INP(n7122), .Z(n7135));
   NBUFFX2 U5897 (.INP(n7121), .Z(n7132));
   NBUFFX2 U5898 (.INP(n7120), .Z(n7131));
   NBUFFX2 U5899 (.INP(n7121), .Z(n7133));
   NBUFFX2 U5900 (.INP(n7119), .Z(n7127));
   NBUFFX2 U5901 (.INP(n7119), .Z(n7126));
   NBUFFX2 U5902 (.INP(n7121), .Z(n7134));
   NBUFFX2 U5903 (.INP(n7120), .Z(n7130));
   NBUFFX2 U5904 (.INP(n7120), .Z(n7129));
   NBUFFX2 U5905 (.INP(n7125), .Z(n7145));
   NBUFFX2 U5906 (.INP(n7125), .Z(n7144));
   NBUFFX2 U5907 (.INP(n7124), .Z(n7143));
   NBUFFX2 U5908 (.INP(n7124), .Z(n7142));
   NBUFFX2 U5909 (.INP(n7124), .Z(n7141));
   NBUFFX2 U5910 (.INP(n7123), .Z(n7140));
   NBUFFX2 U5911 (.INP(n7123), .Z(n7139));
   NBUFFX2 U5912 (.INP(n7123), .Z(n7138));
   NBUFFX2 U5913 (.INP(n7122), .Z(n7137));
   NBUFFX2 U5914 (.INP(n2297), .Z(n7070));
   NBUFFX2 U5915 (.INP(n2298), .Z(n7059));
   NBUFFX2 U5916 (.INP(n7125), .Z(n7146));
   NBUFFX2 U5917 (.INP(n2298), .Z(n7060));
   NBUFFX2 U5918 (.INP(n2298), .Z(n7061));
   NBUFFX2 U5919 (.INP(n2298), .Z(n7062));
   NBUFFX2 U5920 (.INP(n2298), .Z(n7057));
   NBUFFX2 U5921 (.INP(n2298), .Z(n7058));
   NBUFFX2 U5922 (.INP(n7063), .Z(n7038));
   NBUFFX2 U5923 (.INP(n2298), .Z(n7063));
   INVX0 U5924 (.INP(n6966), .ZN(n2276));
   NBUFFX2 U5925 (.INP(n7119), .Z(n7128));
   NOR2X0 U5926 (.IN1(n3410), .IN2(n3411), .QN(n3412));
   NBUFFX2 U5927 (.INP(n7094), .Z(n7108));
   NBUFFX2 U5928 (.INP(n7094), .Z(n7109));
   NBUFFX2 U5929 (.INP(n7095), .Z(n7110));
   NBUFFX2 U5930 (.INP(n7095), .Z(n7111));
   NBUFFX2 U5931 (.INP(n7095), .Z(n7112));
   NBUFFX2 U5932 (.INP(n7096), .Z(n7113));
   NBUFFX2 U5933 (.INP(n7096), .Z(n7114));
   NBUFFX2 U5934 (.INP(n7096), .Z(n7115));
   NBUFFX2 U5935 (.INP(n2297), .Z(n7067));
   NBUFFX2 U5936 (.INP(n2297), .Z(n7066));
   NBUFFX2 U5937 (.INP(n2297), .Z(n7065));
   NBUFFX2 U5938 (.INP(n2297), .Z(n7064));
   NBUFFX2 U5939 (.INP(n7091), .Z(n7098));
   NBUFFX2 U5940 (.INP(n7091), .Z(n7099));
   NBUFFX2 U5941 (.INP(n7091), .Z(n7100));
   NBUFFX2 U5942 (.INP(n7092), .Z(n7101));
   NBUFFX2 U5943 (.INP(n7092), .Z(n7102));
   NBUFFX2 U5944 (.INP(n7092), .Z(n7103));
   NBUFFX2 U5945 (.INP(n7093), .Z(n7104));
   NBUFFX2 U5946 (.INP(n7093), .Z(n7105));
   NBUFFX2 U5947 (.INP(n7093), .Z(n7106));
   NBUFFX2 U5948 (.INP(n7094), .Z(n7107));
   NBUFFX2 U5949 (.INP(n3395), .Z(n6959));
   NBUFFX2 U5950 (.INP(n3395), .Z(n6958));
   NBUFFX2 U5951 (.INP(n3395), .Z(n6957));
   NBUFFX2 U5952 (.INP(n3395), .Z(n6960));
   INVX0 U5953 (.INP(N31), .ZN(n6471));
   INVX0 U5954 (.INP(N30), .ZN(n6472));
   INVX0 U5955 (.INP(N28), .ZN(n6473));
   INVX0 U5956 (.INP(n2966), .ZN(n7583));
   NBUFFX2 U5957 (.INP(n2292), .Z(n7122));
   INVX0 U5958 (.INP(n2941), .ZN(n7581));
   AND2X1 U5959 (.IN1(n3406), .IN2(n3403), .Q(n3401));
   INVX0 U5960 (.INP(n2951), .ZN(n7588));
   NBUFFX2 U5961 (.INP(n2292), .Z(n7121));
   NBUFFX2 U5962 (.INP(n2292), .Z(n7120));
   NBUFFX2 U5963 (.INP(n2292), .Z(n7119));
   INVX0 U5964 (.INP(n2960), .ZN(n7585));
   INVX0 U5965 (.INP(n2963), .ZN(n7584));
   INVX0 U5966 (.INP(n2954), .ZN(n7587));
   NBUFFX2 U5967 (.INP(n2292), .Z(n7125));
   NBUFFX2 U5968 (.INP(n2292), .Z(n7124));
   NBUFFX2 U5969 (.INP(n2292), .Z(n7123));
   OR2X1 U5970 (.IN1(n2941), .IN2(n3403), .Q(n6966));
   INVX0 U5971 (.INP(n3018), .ZN(n7590));
   XOR2X1 U5972 (.IN1(new_sboxw[5]), .IN2(n3072), .Q(n2548));
   XOR2X1 U5973 (.IN1(new_sboxw[1]), .IN2(n3084), .Q(n2568));
   AND3X1 U5974 (.IN1(n3403), .IN2(n7622), .IN3(n7581), .Q(n2298));
   XOR2X1 U5975 (.IN1(new_sboxw[7]), .IN2(n3066), .Q(n2538));
   XOR2X1 U5976 (.IN1(new_sboxw[2]), .IN2(n3081), .Q(n2563));
   XOR2X1 U5977 (.IN1(new_sboxw[5]), .IN2(n3096), .Q(n2586));
   XOR2X1 U5978 (.IN1(new_sboxw[1]), .IN2(n3108), .Q(n2606));
   XOR2X1 U5979 (.IN1(new_sboxw[7]), .IN2(n3090), .Q(n2576));
   XOR2X1 U5980 (.IN1(new_sboxw[2]), .IN2(n3105), .Q(n2601));
   AO21X1 U5981 (.IN1(n7581), .IN2(n7622), .IN3(n2278), .Q(n3405));
   XOR2X1 U5982 (.IN1(new_sboxw[22]), .IN2(n3045), .Q(n2501));
   AND2X1 U5983 (.IN1(n2931), .IN2(n2932), .Q(n6988));
   AND2X1 U5984 (.IN1(n2933), .IN2(n2932), .Q(n6989));
   AND2X1 U5985 (.IN1(n2933), .IN2(n2932), .Q(n6806));
   AND2X1 U5986 (.IN1(n2933), .IN2(n2932), .Q(n6807));
   AND2X1 U5987 (.IN1(n3420), .IN2(n2941), .Q(n3419));
   AO221X1 U5988 (.IN1(n7131), .IN2(n2651), .IN3(key[184]), .IN4(n7309), .IN5(n2652), .Q(
          n2650));
   NOR2X0 U5989 (.IN1(n3397), .IN2(n2214), .QN(n2292));
   AO221X1 U5990 (.IN1(n7136), .IN2(n2926), .IN3(key[129]), .IN4(n7312), .IN5(n2927), .Q(
          n2925));
   AO221X1 U5991 (.IN1(n7136), .IN2(n2901), .IN3(key[134]), .IN4(n2276), .IN5(n2902), .Q(
          n2900));
   AO221X1 U5992 (.IN1(n7136), .IN2(n2911), .IN3(key[132]), .IN4(n7294), .IN5(n2912), .Q(
          n2910));
   NAND2X1 U5993 (.IN1(n3196), .IN2(n3197), .QN(n5431));
   NAND2X1 U5994 (.IN1(n3192), .IN2(n3193), .QN(n5430));
   NAND2X1 U5995 (.IN1(n3188), .IN2(n3189), .QN(n5429));
   NAND2X1 U5996 (.IN1(n3184), .IN2(n3185), .QN(n5428));
   NAND2X1 U5997 (.IN1(n3180), .IN2(n3181), .QN(n5427));
   NAND2X1 U5998 (.IN1(n3132), .IN2(n3133), .QN(n5415));
   NAND2X1 U5999 (.IN1(n3103), .IN2(n3104), .QN(n5407));
   NAND2X1 U6000 (.IN1(n3100), .IN2(n3101), .QN(n5406));
   NAND2X1 U6001 (.IN1(n3097), .IN2(n3098), .QN(n5405));
   NAND2X1 U6002 (.IN1(n3094), .IN2(n3095), .QN(n5404));
   NAND2X1 U6003 (.IN1(n3091), .IN2(n3092), .QN(n5403));
   NAND2X1 U6004 (.IN1(n3073), .IN2(n3074), .QN(n5397));
   NAND2X1 U6005 (.IN1(n3009), .IN2(n3010), .QN(n5375));
   NAND2X1 U6006 (.IN1(n3007), .IN2(n3008), .QN(n5374));
   NAND2X1 U6007 (.IN1(n3005), .IN2(n3006), .QN(n5373));
   NAND2X1 U6008 (.IN1(n3003), .IN2(n3004), .QN(n5372));
   NAND2X1 U6009 (.IN1(n3001), .IN2(n3002), .QN(n5371));
   NAND2X1 U6010 (.IN1(n2999), .IN2(n3000), .QN(n5370));
   NAND2X1 U6011 (.IN1(n2997), .IN2(n2998), .QN(n5369));
   NAND2X1 U6012 (.IN1(n3172), .IN2(n3173), .QN(n5425));
   NAND2X1 U6013 (.IN1(n3168), .IN2(n3169), .QN(n5424));
   NAND2X1 U6014 (.IN1(n3164), .IN2(n3165), .QN(n5423));
   NAND2X1 U6015 (.IN1(n3160), .IN2(n3161), .QN(n5422));
   NAND2X1 U6016 (.IN1(n3156), .IN2(n3157), .QN(n5421));
   NAND2X1 U6017 (.IN1(n3152), .IN2(n3153), .QN(n5420));
   NAND2X1 U6018 (.IN1(n3148), .IN2(n3149), .QN(n5419));
   NAND2X1 U6019 (.IN1(n3144), .IN2(n3145), .QN(n5418));
   NAND2X1 U6020 (.IN1(n3140), .IN2(n3141), .QN(n5417));
   NAND2X1 U6021 (.IN1(n3136), .IN2(n3137), .QN(n5416));
   NAND2X1 U6022 (.IN1(n3128), .IN2(n3129), .QN(n5414));
   NAND2X1 U6023 (.IN1(n3124), .IN2(n3125), .QN(n5413));
   NAND2X1 U6024 (.IN1(n3120), .IN2(n3121), .QN(n5412));
   NAND2X1 U6025 (.IN1(n3116), .IN2(n3117), .QN(n5411));
   NAND2X1 U6026 (.IN1(n3112), .IN2(n3113), .QN(n5410));
   NAND2X1 U6027 (.IN1(n3109), .IN2(n3110), .QN(n5409));
   NAND2X1 U6028 (.IN1(n3106), .IN2(n3107), .QN(n5408));
   NAND2X1 U6029 (.IN1(n3088), .IN2(n3089), .QN(n5402));
   NAND2X1 U6030 (.IN1(n3085), .IN2(n3086), .QN(n5401));
   NAND2X1 U6031 (.IN1(n3082), .IN2(n3083), .QN(n5400));
   NAND2X1 U6032 (.IN1(n3079), .IN2(n3080), .QN(n5399));
   NAND2X1 U6033 (.IN1(n3076), .IN2(n3077), .QN(n5398));
   NAND2X1 U6034 (.IN1(n3067), .IN2(n3068), .QN(n5395));
   NAND2X1 U6035 (.IN1(n3064), .IN2(n3065), .QN(n5394));
   NAND2X1 U6036 (.IN1(n3061), .IN2(n3062), .QN(n5393));
   NAND2X1 U6037 (.IN1(n3058), .IN2(n3059), .QN(n5392));
   NAND2X1 U6038 (.IN1(n3055), .IN2(n3056), .QN(n5391));
   NAND2X1 U6039 (.IN1(n3052), .IN2(n3053), .QN(n5390));
   NAND2X1 U6040 (.IN1(n3049), .IN2(n3050), .QN(n5389));
   NAND2X1 U6041 (.IN1(n3046), .IN2(n3047), .QN(n5388));
   NAND2X1 U6042 (.IN1(n3043), .IN2(n3044), .QN(n5387));
   NAND2X1 U6043 (.IN1(n3040), .IN2(n3041), .QN(n5386));
   NAND2X1 U6044 (.IN1(n3037), .IN2(n3038), .QN(n5385));
   NAND2X1 U6045 (.IN1(n3034), .IN2(n3035), .QN(n5384));
   NAND2X1 U6046 (.IN1(n3031), .IN2(n3032), .QN(n5383));
   NAND2X1 U6047 (.IN1(n3028), .IN2(n3029), .QN(n5382));
   NAND2X1 U6048 (.IN1(n3025), .IN2(n3026), .QN(n5381));
   NAND2X1 U6049 (.IN1(n3022), .IN2(n3023), .QN(n5380));
   NAND2X1 U6050 (.IN1(n3019), .IN2(n3020), .QN(n5379));
   NAND2X1 U6051 (.IN1(n3015), .IN2(n3016), .QN(n5378));
   NAND2X1 U6052 (.IN1(n3013), .IN2(n3014), .QN(n5377));
   NAND2X1 U6053 (.IN1(n3011), .IN2(n3012), .QN(n5376));
   NAND2X1 U6054 (.IN1(n2993), .IN2(n2994), .QN(n5367));
   NAND2X1 U6055 (.IN1(n2991), .IN2(n2992), .QN(n5366));
   NAND2X1 U6056 (.IN1(n2989), .IN2(n2990), .QN(n5365));
   NAND2X1 U6057 (.IN1(n3176), .IN2(n3177), .QN(n5426));
   NAND2X1 U6058 (.IN1(n3070), .IN2(n3071), .QN(n5396));
   NAND2X1 U6059 (.IN1(n2995), .IN2(n2996), .QN(n5368));
   NAND2X1 U6060 (.IN1(n3236), .IN2(n3237), .QN(n5441));
   NAND2X1 U6061 (.IN1(n3232), .IN2(n3233), .QN(n5440));
   NAND2X1 U6062 (.IN1(n3228), .IN2(n3229), .QN(n5439));
   NAND2X1 U6063 (.IN1(n3224), .IN2(n3225), .QN(n5438));
   NAND2X1 U6064 (.IN1(n3220), .IN2(n3221), .QN(n5437));
   NAND2X1 U6065 (.IN1(n3216), .IN2(n3217), .QN(n5436));
   NAND2X1 U6066 (.IN1(n3212), .IN2(n3213), .QN(n5435));
   NAND2X1 U6067 (.IN1(n3270), .IN2(n3271), .QN(n5448));
   NAND2X1 U6068 (.IN1(n3265), .IN2(n3266), .QN(n5447));
   NAND2X1 U6069 (.IN1(n3260), .IN2(n3261), .QN(n5446));
   NAND2X1 U6070 (.IN1(n3255), .IN2(n3256), .QN(n5445));
   NAND2X1 U6071 (.IN1(n3250), .IN2(n3251), .QN(n5444));
   NAND2X1 U6072 (.IN1(n3245), .IN2(n3246), .QN(n5443));
   NAND2X1 U6073 (.IN1(n3240), .IN2(n3241), .QN(n5442));
   NAND2X1 U6074 (.IN1(n3208), .IN2(n3209), .QN(n5434));
   NAND2X1 U6075 (.IN1(n3204), .IN2(n3205), .QN(n5433));
   NAND2X1 U6076 (.IN1(n3200), .IN2(n3201), .QN(n5432));
   AO221X1 U6077 (.IN1(n7131), .IN2(n2626), .IN3(key[189]), .IN4(n7300), .IN5(n2627), .Q(
          n2625));
   AO221X1 U6078 (.IN1(n7135), .IN2(n2886), .IN3(key[137]), .IN4(n7306), .IN5(n2887), .Q(
          n2885));
   AO221X1 U6079 (.IN1(n7132), .IN2(n2681), .IN3(key[178]), .IN4(n7293), .IN5(n2682), .Q(
          n2680));
   AO221X1 U6080 (.IN1(n7135), .IN2(n2841), .IN3(key[146]), .IN4(n7299), .IN5(n2842), .Q(
          n2840));
   AO221X1 U6081 (.IN1(n7133), .IN2(n2741), .IN3(key[166]), .IN4(n7290), .IN5(n2742), .Q(
          n2740));
   AO221X1 U6082 (.IN1(n7133), .IN2(n2721), .IN3(key[170]), .IN4(n2276), .IN5(n2722), .Q(
          n2720));
   AO221X1 U6083 (.IN1(n7135), .IN2(n2866), .IN3(key[141]), .IN4(n2276), .IN5(n2867), .Q(
          n2865));
   AO221X1 U6084 (.IN1(n7133), .IN2(n2726), .IN3(key[169]), .IN4(n7294), .IN5(n2727), .Q(
          n2725));
   AO221X1 U6085 (.IN1(n7131), .IN2(n2646), .IN3(key[185]), .IN4(n7311), .IN5(n2647), .Q(
          n2645));
   AO221X1 U6086 (.IN1(n7135), .IN2(n2881), .IN3(key[138]), .IN4(n7312), .IN5(n2882), .Q(
          n2880));
   AO221X1 U6087 (.IN1(n7133), .IN2(n2766), .IN3(key[161]), .IN4(n7295), .IN5(n2767), .Q(
          n2765));
   AO221X1 U6088 (.IN1(n7131), .IN2(n2631), .IN3(key[188]), .IN4(n7308), .IN5(n2632), .Q(
          n2630));
   AO221X1 U6089 (.IN1(n7131), .IN2(n2641), .IN3(key[186]), .IN4(n7305), .IN5(n2642), .Q(
          n2640));
   AO221X1 U6090 (.IN1(n7127), .IN2(n2406), .IN3(key[233]), .IN4(n7311), .IN5(n2407), .Q(
          n2405));
   AO221X1 U6091 (.IN1(n7126), .IN2(n2341), .IN3(key[246]), .IN4(n7311), .IN5(n2342), .Q(
          n2340));
   AO221X1 U6092 (.IN1(n7127), .IN2(n2401), .IN3(key[234]), .IN4(n7311), .IN5(n2402), .Q(
          n2400));
   AO221X1 U6093 (.IN1(n7126), .IN2(n2311), .IN3(key[252]), .IN4(n7307), .IN5(n2312), .Q(
          n2310));
   AO221X1 U6094 (.IN1(n7126), .IN2(n2306), .IN3(key[253]), .IN4(n7308), .IN5(n2307), .Q(
          n2305));
   AO221X1 U6095 (.IN1(n7126), .IN2(n2293), .IN3(key[255]), .IN4(n7300), .IN5(n2294), .Q(
          n2277));
   AO221X1 U6096 (.IN1(n7127), .IN2(n2361), .IN3(key[242]), .IN4(n7290), .IN5(n2362), .Q(
          n2360));
   AO221X1 U6097 (.IN1(n7127), .IN2(n2411), .IN3(key[232]), .IN4(n7295), .IN5(n2412), .Q(
          n2410));
   AO221X1 U6098 (.IN1(n7127), .IN2(n2396), .IN3(key[235]), .IN4(n7305), .IN5(n2397), .Q(
          n2395));
   AO221X1 U6099 (.IN1(n7127), .IN2(n2386), .IN3(key[237]), .IN4(n7299), .IN5(n2387), .Q(
          n2385));
   AO221X1 U6100 (.IN1(n7128), .IN2(n2451), .IN3(key[224]), .IN4(n7296), .IN5(n2452), .Q(
          n2450));
   XNOR3X1 U6101 (.IN1(n4), .IN2(n7583), .IN3(n2196), .Q(n2814));
   XOR3X1 U6102 (.IN1(sboxw[24]), .IN2(prev_key1_reg[88]), .IN3(prev_key1_reg[56]), .Q(
          n2196));
   AO221X1 U6103 (.IN1(n7128), .IN2(n2446), .IN3(key[225]), .IN4(n7301), .IN5(n2447), .Q(
          n2445));
   NAND2X1 U6104 (.IN1(n2955), .IN2(n2956), .QN(n5350));
   NAND2X1 U6105 (.IN1(n2952), .IN2(n2953), .QN(n5349));
   NAND2X1 U6106 (.IN1(n2949), .IN2(n2950), .QN(n5348));
   NAND2X1 U6107 (.IN1(n2946), .IN2(n2947), .QN(n5347));
   NAND2X1 U6108 (.IN1(n2942), .IN2(n2943), .QN(n5346));
   NAND2X1 U6109 (.IN1(n3365), .IN2(n3366), .QN(n5467));
   NAND2X1 U6110 (.IN1(n3360), .IN2(n3361), .QN(n5466));
   NAND2X1 U6111 (.IN1(n3355), .IN2(n3356), .QN(n5465));
   NAND2X1 U6112 (.IN1(n3350), .IN2(n3351), .QN(n5464));
   NAND2X1 U6113 (.IN1(n3345), .IN2(n3346), .QN(n5463));
   NAND2X1 U6114 (.IN1(n3340), .IN2(n3341), .QN(n5462));
   NAND2X1 U6115 (.IN1(n3335), .IN2(n3336), .QN(n5461));
   NAND2X1 U6116 (.IN1(n3330), .IN2(n3331), .QN(n5460));
   NAND2X1 U6117 (.IN1(n3325), .IN2(n3326), .QN(n5459));
   NAND2X1 U6118 (.IN1(n3320), .IN2(n3321), .QN(n5458));
   NAND2X1 U6119 (.IN1(n3315), .IN2(n3316), .QN(n5457));
   NAND2X1 U6120 (.IN1(n3310), .IN2(n3311), .QN(n5456));
   NAND2X1 U6121 (.IN1(n3305), .IN2(n3306), .QN(n5455));
   NAND2X1 U6122 (.IN1(n3300), .IN2(n3301), .QN(n5454));
   NAND2X1 U6123 (.IN1(n3295), .IN2(n3296), .QN(n5453));
   NAND2X1 U6124 (.IN1(n3290), .IN2(n3291), .QN(n5452));
   NAND2X1 U6125 (.IN1(n3285), .IN2(n3286), .QN(n5451));
   NAND2X1 U6126 (.IN1(n3280), .IN2(n3281), .QN(n5450));
   NAND2X1 U6127 (.IN1(n3275), .IN2(n3276), .QN(n5449));
   NAND2X1 U6128 (.IN1(n2987), .IN2(n2988), .QN(n5364));
   NAND2X1 U6129 (.IN1(n2985), .IN2(n2986), .QN(n5363));
   NAND2X1 U6130 (.IN1(n2983), .IN2(n2984), .QN(n5362));
   NAND2X1 U6131 (.IN1(n2981), .IN2(n2982), .QN(n5361));
   NAND2X1 U6132 (.IN1(n2979), .IN2(n2980), .QN(n5360));
   NAND2X1 U6133 (.IN1(n2977), .IN2(n2978), .QN(n5359));
   NAND2X1 U6134 (.IN1(n2975), .IN2(n2976), .QN(n5358));
   NAND2X1 U6135 (.IN1(n2973), .IN2(n2974), .QN(n5357));
   NAND2X1 U6136 (.IN1(n2971), .IN2(n2972), .QN(n5356));
   NAND2X1 U6137 (.IN1(n2969), .IN2(n2970), .QN(n5355));
   NAND2X1 U6138 (.IN1(n2967), .IN2(n2968), .QN(n5354));
   NAND2X1 U6139 (.IN1(n2964), .IN2(n2965), .QN(n5353));
   NAND2X1 U6140 (.IN1(n2961), .IN2(n2962), .QN(n5352));
   NAND2X1 U6141 (.IN1(n2958), .IN2(n2959), .QN(n5351));
   XNOR3X1 U6142 (.IN1(n2198), .IN2(new_sboxw[5]), .IN3(n2197), .Q(n2709));
   XOR2X1 U6143 (.IN1(prev_key1_reg[45]), .IN2(prev_key1_reg[77]), .Q(n2197));
   XNOR3X1 U6144 (.IN1(n2198), .IN2(new_sboxw[5]), .IN3(n2199), .Q(n2869));
   XOR3X1 U6145 (.IN1(sboxw[13]), .IN2(prev_key1_reg[77]), .IN3(prev_key1_reg[45]), .Q(
          n2199));
   XNOR3X1 U6146 (.IN1(n2200), .IN2(new_sboxw[7]), .IN3(n2201), .Q(n2859));
   XOR3X1 U6147 (.IN1(sboxw[15]), .IN2(prev_key1_reg[79]), .IN3(prev_key1_reg[47]), .Q(
          n2201));
   XNOR3X1 U6148 (.IN1(n2202), .IN2(new_sboxw[2]), .IN3(n2203), .Q(n2884));
   XOR3X1 U6149 (.IN1(sboxw[10]), .IN2(prev_key1_reg[74]), .IN3(prev_key1_reg[42]), .Q(
          n2203));
   XOR3X1 U6150 (.IN1(prev_key1_reg[77]), .IN2(prev_key1_reg[109]), .IN3(new_sboxw[5]), .Q(
          n2549));
   XOR3X1 U6151 (.IN1(prev_key1_reg[73]), .IN2(prev_key1_reg[105]), .IN3(new_sboxw[1]), .Q(
          n2569));
   NAND2X1 U6152 (.IN1(n3398), .IN2(n3399), .QN(n5601));
   NAND2X1 U6153 (.IN1(n3390), .IN2(n3391), .QN(n5472));
   NAND2X1 U6154 (.IN1(n3385), .IN2(n3386), .QN(n5471));
   NAND2X1 U6155 (.IN1(n3380), .IN2(n3381), .QN(n5470));
   NAND2X1 U6156 (.IN1(n3375), .IN2(n3376), .QN(n5469));
   NAND2X1 U6157 (.IN1(n3370), .IN2(n3371), .QN(n5468));
   XOR3X1 U6158 (.IN1(prev_key1_reg[79]), .IN2(prev_key1_reg[111]), .IN3(new_sboxw[7]), .Q(
          n2539));
   XOR3X1 U6159 (.IN1(prev_key1_reg[74]), .IN2(prev_key1_reg[106]), .IN3(new_sboxw[2]), .Q(
          n2564));
   XNOR2X1 U6160 (.IN1(new_sboxw[22]), .IN2(n2224), .Q(n2341));
   NAND3X0 U6161 (.IN1(n2934), .IN2(n2933), .IN3(round_ctr_reg[3]), .QN(n2290));
   NAND3X0 U6162 (.IN1(n2933), .IN2(n2212), .IN3(n2934), .QN(n2282));
   NAND3X0 U6163 (.IN1(n2933), .IN2(round_ctr_reg[1]), .IN3(n2936), .QN(n2288));
   NAND3X0 U6164 (.IN1(n2933), .IN2(n2213), .IN3(n2936), .QN(n2286));
   AND4X1 U6165 (.IN1(round_ctr_reg[3]), .IN2(round_ctr_reg[2]), .IN3(n2931), .IN4(
          round_ctr_reg[1]), .Q(n6992));
   AND2X1 U6166 (.IN1(round_ctr_reg[2]), .IN2(n2213), .Q(n2934));
   NAND3X0 U6167 (.IN1(n2934), .IN2(n2931), .IN3(round_ctr_reg[3]), .QN(n2289));
   AND3X1 U6168 (.IN1(n2931), .IN2(round_ctr_reg[1]), .IN3(n2936), .Q(n6991));
   AND3X1 U6169 (.IN1(n2931), .IN2(n2213), .IN3(n2936), .Q(n6993));
   XNOR2X1 U6170 (.IN1(keylen), .IN2(round_ctr_reg[2]), .Q(n3425));
   AOI221X1 U6171 (.IN1(n3423), .IN2(key_mem_ctrl_reg[1]), .IN3(init), .IN4(n2242), .IN5(
          key_mem_ctrl_reg[0]), .QN(n2204));
   NAND3X0 U6172 (.IN1(n3420), .IN2(n2941), .IN3(n3421), .QN(n5615));
   NAND2X0 U6173 (.IN1(key_mem_ctrl_reg[1]), .IN2(n2204), .QN(n3421));
   INVX0 U6174 (.INP(n3408), .ZN(n7582));
   NAND2X1 U6175 (.IN1(n2242), .IN2(key_mem_ctrl_reg[0]), .QN(n3420));
   NOR2X0 U6176 (.IN1(n6472), .IN2(N31), .QN(n2231));
   NOR2X0 U6177 (.IN1(N28), .IN2(N29), .QN(n2209));
   AND2X1 U6178 (.IN1(n2231), .IN2(n2209), .Q(n6453));
   NOR2X0 U6179 (.IN1(n6473), .IN2(N29), .QN(n2210));
   AND2X1 U6180 (.IN1(n2231), .IN2(n2210), .Q(n6452));
   AND2X1 U6181 (.IN1(N28), .IN2(N29), .Q(n2211));
   NOR2X0 U6182 (.IN1(n6471), .IN2(N30), .QN(n2206));
   AND2X1 U6183 (.IN1(n2211), .IN2(n2206), .Q(n6450));
   AND2X1 U6184 (.IN1(N29), .IN2(n6473), .Q(n2232));
   AND2X1 U6185 (.IN1(n2231), .IN2(n2232), .Q(n6449));
   AO22X1 U6186 (.IN1(\key_mem[11][0] ), .IN2(n6499), .IN3(\key_mem[6][0] ), .IN4(n6484), .
          Q(n2205));
   AO221X1 U6187 (.IN1(\key_mem[4][0] ), .IN2(n6529), .IN3(\key_mem[5][0] ), .IN4(n6514), .
          IN5(n2205), .Q(n2238));
   AND2X1 U6188 (.IN1(n2210), .IN2(n2206), .Q(n6456));
   AND2X1 U6189 (.IN1(n2209), .IN2(n2206), .Q(n6455));
   AND2X1 U6190 (.IN1(n2206), .IN2(n2232), .Q(n6454));
   AO222X1 U6191 (.IN1(\key_mem[9][0] ), .IN2(n6574), .IN3(\key_mem[8][0] ), .IN4(n6559), .
          IN5(\key_mem[10][0] ), .IN6(n6544), .Q(n2237));
   NOR2X0 U6192 (.IN1(n6472), .IN2(n6471), .QN(n2207));
   AND2X1 U6193 (.IN1(n2207), .IN2(n2209), .Q(n6461));
   AND2X1 U6194 (.IN1(n2207), .IN2(n2210), .Q(n6460));
   NOR2X0 U6195 (.IN1(N30), .IN2(N31), .QN(n2233));
   AND2X1 U6196 (.IN1(n2233), .IN2(n2211), .Q(n6458));
   AND2X1 U6197 (.IN1(n2207), .IN2(n2232), .Q(n6457));
   AO22X1 U6198 (.IN1(\key_mem[3][0] ), .IN2(n6604), .IN3(\key_mem[14][0] ), .IN4(n6589), .
          Q(n2208));
   AO221X1 U6199 (.IN1(\key_mem[12][0] ), .IN2(n6634), .IN3(\key_mem[13][0] ), .IN4(n6619)
          , .IN5(n2208), .Q(n2236));
   AND2X1 U6200 (.IN1(n2233), .IN2(n2209), .Q(n6466));
   AND2X1 U6201 (.IN1(n2233), .IN2(n2210), .Q(n6465));
   AND2X1 U6202 (.IN1(n2231), .IN2(n2211), .Q(n6463));
   AO22X1 U6203 (.IN1(\key_mem[7][0] ), .IN2(n6664), .IN3(\key_mem[2][0] ), .IN4(n6649), .
          Q(n2234));
   AO221X1 U6204 (.IN1(\key_mem[0][0] ), .IN2(n6694), .IN3(\key_mem[1][0] ), .IN4(n6679), .
          IN5(n2234), .Q(n2235));
   OR4X1 U6205 (.IN1(n2238), .IN2(n2237), .IN3(n2236), .IN4(n2235), .Q(round_key[0]));
   AO22X1 U6206 (.IN1(\key_mem[11][1] ), .IN2(n6499), .IN3(\key_mem[6][1] ), .IN4(n6484), .
          Q(n2239));
   AO221X1 U6207 (.IN1(\key_mem[4][1] ), .IN2(n6529), .IN3(\key_mem[5][1] ), .IN4(n6514), .
          IN5(n2239), .Q(n2247));
   AO222X1 U6208 (.IN1(\key_mem[9][1] ), .IN2(n6574), .IN3(\key_mem[8][1] ), .IN4(n6559), .
          IN5(\key_mem[10][1] ), .IN6(n6544), .Q(n2246));
   AO22X1 U6209 (.IN1(\key_mem[3][1] ), .IN2(n6604), .IN3(\key_mem[14][1] ), .IN4(n6589), .
          Q(n2240));
   AO221X1 U6210 (.IN1(\key_mem[12][1] ), .IN2(n6634), .IN3(\key_mem[13][1] ), .IN4(n6619)
          , .IN5(n2240), .Q(n2245));
   AO22X1 U6211 (.IN1(\key_mem[7][1] ), .IN2(n6664), .IN3(\key_mem[2][1] ), .IN4(n6649), .
          Q(n2241));
   AO221X1 U6212 (.IN1(\key_mem[0][1] ), .IN2(n6694), .IN3(\key_mem[1][1] ), .IN4(n6679), .
          IN5(n2241), .Q(n2244));
   OR4X1 U6213 (.IN1(n2247), .IN2(n2246), .IN3(n2245), .IN4(n2244), .Q(round_key[1]));
   AO22X1 U6214 (.IN1(\key_mem[11][2] ), .IN2(n6499), .IN3(\key_mem[6][2] ), .IN4(n6484), .
          Q(n2248));
   AO221X1 U6215 (.IN1(\key_mem[4][2] ), .IN2(n6529), .IN3(\key_mem[5][2] ), .IN4(n6514), .
          IN5(n2248), .Q(n2254));
   AO222X1 U6216 (.IN1(\key_mem[9][2] ), .IN2(n6574), .IN3(\key_mem[8][2] ), .IN4(n6559), .
          IN5(\key_mem[10][2] ), .IN6(n6544), .Q(n2253));
   AO22X1 U6217 (.IN1(\key_mem[3][2] ), .IN2(n6604), .IN3(\key_mem[14][2] ), .IN4(n6589), .
          Q(n2249));
   AO221X1 U6218 (.IN1(\key_mem[12][2] ), .IN2(n6634), .IN3(\key_mem[13][2] ), .IN4(n6619)
          , .IN5(n2249), .Q(n2252));
   AO22X1 U6219 (.IN1(\key_mem[7][2] ), .IN2(n6664), .IN3(\key_mem[2][2] ), .IN4(n6649), .
          Q(n2250));
   AO221X1 U6220 (.IN1(\key_mem[0][2] ), .IN2(n6694), .IN3(\key_mem[1][2] ), .IN4(n6679), .
          IN5(n2250), .Q(n2251));
   OR4X1 U6221 (.IN1(n2254), .IN2(n2253), .IN3(n2252), .IN4(n2251), .Q(round_key[2]));
   AO22X1 U6222 (.IN1(\key_mem[11][3] ), .IN2(n6499), .IN3(\key_mem[6][3] ), .IN4(n6484), .
          Q(n2255));
   AO221X1 U6223 (.IN1(\key_mem[4][3] ), .IN2(n6529), .IN3(\key_mem[5][3] ), .IN4(n6514), .
          IN5(n2255), .Q(n2261));
   AO222X1 U6224 (.IN1(\key_mem[9][3] ), .IN2(n6574), .IN3(\key_mem[8][3] ), .IN4(n6559), .
          IN5(\key_mem[10][3] ), .IN6(n6544), .Q(n2260));
   AO22X1 U6225 (.IN1(\key_mem[3][3] ), .IN2(n6604), .IN3(\key_mem[14][3] ), .IN4(n6589), .
          Q(n2256));
   AO221X1 U6226 (.IN1(\key_mem[12][3] ), .IN2(n6634), .IN3(\key_mem[13][3] ), .IN4(n6619)
          , .IN5(n2256), .Q(n2259));
   AO22X1 U6227 (.IN1(\key_mem[7][3] ), .IN2(n6664), .IN3(\key_mem[2][3] ), .IN4(n6649), .
          Q(n2257));
   AO221X1 U6228 (.IN1(\key_mem[0][3] ), .IN2(n6694), .IN3(\key_mem[1][3] ), .IN4(n6679), .
          IN5(n2257), .Q(n2258));
   OR4X1 U6229 (.IN1(n2261), .IN2(n2260), .IN3(n2259), .IN4(n2258), .Q(round_key[3]));
   AO22X1 U6230 (.IN1(\key_mem[11][4] ), .IN2(n6499), .IN3(\key_mem[6][4] ), .IN4(n6484), .
          Q(n2262));
   AO221X1 U6231 (.IN1(\key_mem[4][4] ), .IN2(n6529), .IN3(\key_mem[5][4] ), .IN4(n6514), .
          IN5(n2262), .Q(n2268));
   AO222X1 U6232 (.IN1(\key_mem[9][4] ), .IN2(n6574), .IN3(\key_mem[8][4] ), .IN4(n6559), .
          IN5(\key_mem[10][4] ), .IN6(n6544), .Q(n2267));
   AO22X1 U6233 (.IN1(\key_mem[3][4] ), .IN2(n6604), .IN3(\key_mem[14][4] ), .IN4(n6589), .
          Q(n2263));
   AO221X1 U6234 (.IN1(\key_mem[12][4] ), .IN2(n6634), .IN3(\key_mem[13][4] ), .IN4(n6619)
          , .IN5(n2263), .Q(n2266));
   AO22X1 U6235 (.IN1(\key_mem[7][4] ), .IN2(n6664), .IN3(\key_mem[2][4] ), .IN4(n6649), .
          Q(n2264));
   AO221X1 U6236 (.IN1(\key_mem[0][4] ), .IN2(n6694), .IN3(\key_mem[1][4] ), .IN4(n6679), .
          IN5(n2264), .Q(n2265));
   OR4X1 U6237 (.IN1(n2268), .IN2(n2267), .IN3(n2266), .IN4(n2265), .Q(round_key[4]));
   AO22X1 U6238 (.IN1(\key_mem[11][5] ), .IN2(n6499), .IN3(\key_mem[6][5] ), .IN4(n6484), .
          Q(n2269));
   AO221X1 U6239 (.IN1(\key_mem[4][5] ), .IN2(n6529), .IN3(\key_mem[5][5] ), .IN4(n6514), .
          IN5(n2269), .Q(n2275));
   AO222X1 U6240 (.IN1(\key_mem[9][5] ), .IN2(n6574), .IN3(\key_mem[8][5] ), .IN4(n6559), .
          IN5(\key_mem[10][5] ), .IN6(n6544), .Q(n2274));
   AO22X1 U6241 (.IN1(\key_mem[3][5] ), .IN2(n6604), .IN3(\key_mem[14][5] ), .IN4(n6589), .
          Q(n2270));
   AO221X1 U6242 (.IN1(\key_mem[12][5] ), .IN2(n6634), .IN3(\key_mem[13][5] ), .IN4(n6619)
          , .IN5(n2270), .Q(n2273));
   AO22X1 U6243 (.IN1(\key_mem[7][5] ), .IN2(n6664), .IN3(\key_mem[2][5] ), .IN4(n6649), .
          Q(n2271));
   AO221X1 U6244 (.IN1(\key_mem[0][5] ), .IN2(n6694), .IN3(\key_mem[1][5] ), .IN4(n6679), .
          IN5(n2271), .Q(n2272));
   OR4X1 U6245 (.IN1(n2275), .IN2(n2274), .IN3(n2273), .IN4(n2272), .Q(round_key[5]));
   AO22X1 U6246 (.IN1(\key_mem[11][6] ), .IN2(n6499), .IN3(\key_mem[6][6] ), .IN4(n6484), .
          Q(n2279));
   AO221X1 U6247 (.IN1(\key_mem[4][6] ), .IN2(n6529), .IN3(\key_mem[5][6] ), .IN4(n6514), .
          IN5(n2279), .Q(n3143));
   AO222X1 U6248 (.IN1(\key_mem[9][6] ), .IN2(n6574), .IN3(\key_mem[8][6] ), .IN4(n6559), .
          IN5(\key_mem[10][6] ), .IN6(n6544), .Q(n2291));
   AO22X1 U6249 (.IN1(\key_mem[3][6] ), .IN2(n6604), .IN3(\key_mem[14][6] ), .IN4(n6589), .
          Q(n2280));
   AO221X1 U6250 (.IN1(\key_mem[12][6] ), .IN2(n6634), .IN3(\key_mem[13][6] ), .IN4(n6619)
          , .IN5(n2280), .Q(n2287));
   AO22X1 U6251 (.IN1(\key_mem[7][6] ), .IN2(n6664), .IN3(\key_mem[2][6] ), .IN4(n6649), .
          Q(n2281));
   AO221X1 U6252 (.IN1(\key_mem[0][6] ), .IN2(n6694), .IN3(\key_mem[1][6] ), .IN4(n6679), .
          IN5(n2281), .Q(n2285));
   OR4X1 U6253 (.IN1(n3143), .IN2(n2291), .IN3(n2287), .IN4(n2285), .Q(round_key[6]));
   AO22X1 U6254 (.IN1(\key_mem[11][7] ), .IN2(n6499), .IN3(\key_mem[6][7] ), .IN4(n6484), .
          Q(n3187));
   AO221X1 U6255 (.IN1(\key_mem[4][7] ), .IN2(n6529), .IN3(\key_mem[5][7] ), .IN4(n6514), .
          IN5(n3187), .Q(n3422));
   AO222X1 U6256 (.IN1(\key_mem[9][7] ), .IN2(n6574), .IN3(\key_mem[8][7] ), .IN4(n6559), .
          IN5(\key_mem[10][7] ), .IN6(n6544), .Q(n3409));
   AO22X1 U6257 (.IN1(\key_mem[3][7] ), .IN2(n6604), .IN3(\key_mem[14][7] ), .IN4(n6589), .
          Q(n3279));
   AO221X1 U6258 (.IN1(\key_mem[12][7] ), .IN2(n6634), .IN3(\key_mem[13][7] ), .IN4(n6619)
          , .IN5(n3279), .Q(n3349));
   AO22X1 U6259 (.IN1(\key_mem[7][7] ), .IN2(n6664), .IN3(\key_mem[2][7] ), .IN4(n6649), .
          Q(n3324));
   AO221X1 U6260 (.IN1(\key_mem[0][7] ), .IN2(n6694), .IN3(\key_mem[1][7] ), .IN4(n6679), .
          IN5(n3324), .Q(n3334));
   OR4X1 U6261 (.IN1(n3422), .IN2(n3409), .IN3(n3349), .IN4(n3334), .Q(round_key[7]));
   AO22X1 U6262 (.IN1(\key_mem[11][8] ), .IN2(n6499), .IN3(\key_mem[6][8] ), .IN4(n6484), .
          Q(n3424));
   AO221X1 U6263 (.IN1(\key_mem[4][8] ), .IN2(n6529), .IN3(\key_mem[5][8] ), .IN4(n6514), .
          IN5(n3424), .Q(n5622));
   AO222X1 U6264 (.IN1(\key_mem[9][8] ), .IN2(n6574), .IN3(\key_mem[8][8] ), .IN4(n6559), .
          IN5(\key_mem[10][8] ), .IN6(n6544), .Q(n5621));
   AO22X1 U6265 (.IN1(\key_mem[3][8] ), .IN2(n6604), .IN3(\key_mem[14][8] ), .IN4(n6589), .
          Q(n5617));
   AO221X1 U6266 (.IN1(\key_mem[12][8] ), .IN2(n6634), .IN3(\key_mem[13][8] ), .IN4(n6619)
          , .IN5(n5617), .Q(n5620));
   AO22X1 U6267 (.IN1(\key_mem[7][8] ), .IN2(n6664), .IN3(\key_mem[2][8] ), .IN4(n6649), .
          Q(n5618));
   AO221X1 U6268 (.IN1(\key_mem[0][8] ), .IN2(n6694), .IN3(\key_mem[1][8] ), .IN4(n6679), .
          IN5(n5618), .Q(n5619));
   OR4X1 U6269 (.IN1(n5622), .IN2(n5621), .IN3(n5620), .IN4(n5619), .Q(round_key[8]));
   AO22X1 U6270 (.IN1(\key_mem[11][9] ), .IN2(n6499), .IN3(\key_mem[6][9] ), .IN4(n6484), .
          Q(n5623));
   AO221X1 U6271 (.IN1(\key_mem[4][9] ), .IN2(n6529), .IN3(\key_mem[5][9] ), .IN4(n6514), .
          IN5(n5623), .Q(n5629));
   AO222X1 U6272 (.IN1(\key_mem[9][9] ), .IN2(n6574), .IN3(\key_mem[8][9] ), .IN4(n6559), .
          IN5(\key_mem[10][9] ), .IN6(n6544), .Q(n5628));
   AO22X1 U6273 (.IN1(\key_mem[3][9] ), .IN2(n6604), .IN3(\key_mem[14][9] ), .IN4(n6589), .
          Q(n5624));
   AO221X1 U6274 (.IN1(\key_mem[12][9] ), .IN2(n6634), .IN3(\key_mem[13][9] ), .IN4(n6619)
          , .IN5(n5624), .Q(n5627));
   AO22X1 U6275 (.IN1(\key_mem[7][9] ), .IN2(n6664), .IN3(\key_mem[2][9] ), .IN4(n6649), .
          Q(n5625));
   AO221X1 U6276 (.IN1(\key_mem[0][9] ), .IN2(n6694), .IN3(\key_mem[1][9] ), .IN4(n6679), .
          IN5(n5625), .Q(n5626));
   OR4X1 U6277 (.IN1(n5629), .IN2(n5628), .IN3(n5627), .IN4(n5626), .Q(round_key[9]));
   AO22X1 U6278 (.IN1(\key_mem[11][10] ), .IN2(n6499), .IN3(\key_mem[6][10] ), .IN4(n6484)
          , .Q(n5630));
   AO221X1 U6279 (.IN1(\key_mem[4][10] ), .IN2(n6529), .IN3(\key_mem[5][10] ), .IN4(n6514)
          , .IN5(n5630), .Q(n5636));
   AO222X1 U6280 (.IN1(\key_mem[9][10] ), .IN2(n6574), .IN3(\key_mem[8][10] ), .IN4(n6559)
          , .IN5(\key_mem[10][10] ), .IN6(n6544), .Q(n5635));
   AO22X1 U6281 (.IN1(\key_mem[3][10] ), .IN2(n6604), .IN3(\key_mem[14][10] ), .IN4(n6589)
          , .Q(n5631));
   AO221X1 U6282 (.IN1(\key_mem[12][10] ), .IN2(n6634), .IN3(\key_mem[13][10] ), .IN4(
          n6619), .IN5(n5631), .Q(n5634));
   AO22X1 U6283 (.IN1(\key_mem[7][10] ), .IN2(n6664), .IN3(\key_mem[2][10] ), .IN4(n6649)
          , .Q(n5632));
   AO221X1 U6284 (.IN1(\key_mem[0][10] ), .IN2(n6694), .IN3(\key_mem[1][10] ), .IN4(n6679)
          , .IN5(n5632), .Q(n5633));
   OR4X1 U6285 (.IN1(n5636), .IN2(n5635), .IN3(n5634), .IN4(n5633), .Q(round_key[10]));
   AO22X1 U6286 (.IN1(\key_mem[11][11] ), .IN2(n6499), .IN3(\key_mem[6][11] ), .IN4(n6484)
          , .Q(n5637));
   AO221X1 U6287 (.IN1(\key_mem[4][11] ), .IN2(n6529), .IN3(\key_mem[5][11] ), .IN4(n6514)
          , .IN5(n5637), .Q(n5643));
   AO222X1 U6288 (.IN1(\key_mem[9][11] ), .IN2(n6574), .IN3(\key_mem[8][11] ), .IN4(n6559)
          , .IN5(\key_mem[10][11] ), .IN6(n6544), .Q(n5642));
   AO22X1 U6289 (.IN1(\key_mem[3][11] ), .IN2(n6604), .IN3(\key_mem[14][11] ), .IN4(n6589)
          , .Q(n5638));
   AO221X1 U6290 (.IN1(\key_mem[12][11] ), .IN2(n6634), .IN3(\key_mem[13][11] ), .IN4(
          n6619), .IN5(n5638), .Q(n5641));
   AO22X1 U6291 (.IN1(\key_mem[7][11] ), .IN2(n6664), .IN3(\key_mem[2][11] ), .IN4(n6649)
          , .Q(n5639));
   AO221X1 U6292 (.IN1(\key_mem[0][11] ), .IN2(n6694), .IN3(\key_mem[1][11] ), .IN4(n6679)
          , .IN5(n5639), .Q(n5640));
   OR4X1 U6293 (.IN1(n5643), .IN2(n5642), .IN3(n5641), .IN4(n5640), .Q(round_key[11]));
   AO22X1 U6294 (.IN1(\key_mem[11][12] ), .IN2(n6498), .IN3(\key_mem[6][12] ), .IN4(n6483)
          , .Q(n5644));
   AO221X1 U6295 (.IN1(\key_mem[4][12] ), .IN2(n6528), .IN3(\key_mem[5][12] ), .IN4(n6513)
          , .IN5(n5644), .Q(n5650));
   AO222X1 U6296 (.IN1(\key_mem[9][12] ), .IN2(n6573), .IN3(\key_mem[8][12] ), .IN4(n6558)
          , .IN5(\key_mem[10][12] ), .IN6(n6543), .Q(n5649));
   AO22X1 U6297 (.IN1(\key_mem[3][12] ), .IN2(n6603), .IN3(\key_mem[14][12] ), .IN4(n6588)
          , .Q(n5645));
   AO221X1 U6298 (.IN1(\key_mem[12][12] ), .IN2(n6633), .IN3(\key_mem[13][12] ), .IN4(
          n6618), .IN5(n5645), .Q(n5648));
   AO22X1 U6299 (.IN1(\key_mem[7][12] ), .IN2(n6663), .IN3(\key_mem[2][12] ), .IN4(n6648)
          , .Q(n5646));
   AO221X1 U6300 (.IN1(\key_mem[0][12] ), .IN2(n6693), .IN3(\key_mem[1][12] ), .IN4(n6678)
          , .IN5(n5646), .Q(n5647));
   OR4X1 U6301 (.IN1(n5650), .IN2(n5649), .IN3(n5648), .IN4(n5647), .Q(round_key[12]));
   AO22X1 U6302 (.IN1(\key_mem[11][13] ), .IN2(n6498), .IN3(\key_mem[6][13] ), .IN4(n6483)
          , .Q(n5651));
   AO221X1 U6303 (.IN1(\key_mem[4][13] ), .IN2(n6528), .IN3(\key_mem[5][13] ), .IN4(n6513)
          , .IN5(n5651), .Q(n5657));
   AO222X1 U6304 (.IN1(\key_mem[9][13] ), .IN2(n6573), .IN3(\key_mem[8][13] ), .IN4(n6558)
          , .IN5(\key_mem[10][13] ), .IN6(n6543), .Q(n5656));
   AO22X1 U6305 (.IN1(\key_mem[3][13] ), .IN2(n6603), .IN3(\key_mem[14][13] ), .IN4(n6588)
          , .Q(n5652));
   AO221X1 U6306 (.IN1(\key_mem[12][13] ), .IN2(n6633), .IN3(\key_mem[13][13] ), .IN4(
          n6618), .IN5(n5652), .Q(n5655));
   AO22X1 U6307 (.IN1(\key_mem[7][13] ), .IN2(n6663), .IN3(\key_mem[2][13] ), .IN4(n6648)
          , .Q(n5653));
   AO221X1 U6308 (.IN1(\key_mem[0][13] ), .IN2(n6693), .IN3(\key_mem[1][13] ), .IN4(n6678)
          , .IN5(n5653), .Q(n5654));
   OR4X1 U6309 (.IN1(n5657), .IN2(n5656), .IN3(n5655), .IN4(n5654), .Q(round_key[13]));
   AO22X1 U6310 (.IN1(\key_mem[11][14] ), .IN2(n6498), .IN3(\key_mem[6][14] ), .IN4(n6483)
          , .Q(n5658));
   AO221X1 U6311 (.IN1(\key_mem[4][14] ), .IN2(n6528), .IN3(\key_mem[5][14] ), .IN4(n6513)
          , .IN5(n5658), .Q(n5664));
   AO222X1 U6312 (.IN1(\key_mem[9][14] ), .IN2(n6573), .IN3(\key_mem[8][14] ), .IN4(n6558)
          , .IN5(\key_mem[10][14] ), .IN6(n6543), .Q(n5663));
   AO22X1 U6313 (.IN1(\key_mem[3][14] ), .IN2(n6603), .IN3(\key_mem[14][14] ), .IN4(n6588)
          , .Q(n5659));
   AO221X1 U6314 (.IN1(\key_mem[12][14] ), .IN2(n6633), .IN3(\key_mem[13][14] ), .IN4(
          n6618), .IN5(n5659), .Q(n5662));
   AO22X1 U6315 (.IN1(\key_mem[7][14] ), .IN2(n6663), .IN3(\key_mem[2][14] ), .IN4(n6648)
          , .Q(n5660));
   AO221X1 U6316 (.IN1(\key_mem[0][14] ), .IN2(n6693), .IN3(\key_mem[1][14] ), .IN4(n6678)
          , .IN5(n5660), .Q(n5661));
   OR4X1 U6317 (.IN1(n5664), .IN2(n5663), .IN3(n5662), .IN4(n5661), .Q(round_key[14]));
   AO22X1 U6318 (.IN1(\key_mem[11][15] ), .IN2(n6498), .IN3(\key_mem[6][15] ), .IN4(n6483)
          , .Q(n5665));
   AO221X1 U6319 (.IN1(\key_mem[4][15] ), .IN2(n6528), .IN3(\key_mem[5][15] ), .IN4(n6513)
          , .IN5(n5665), .Q(n5671));
   AO222X1 U6320 (.IN1(\key_mem[9][15] ), .IN2(n6573), .IN3(\key_mem[8][15] ), .IN4(n6558)
          , .IN5(\key_mem[10][15] ), .IN6(n6543), .Q(n5670));
   AO22X1 U6321 (.IN1(\key_mem[3][15] ), .IN2(n6603), .IN3(\key_mem[14][15] ), .IN4(n6588)
          , .Q(n5666));
   AO221X1 U6322 (.IN1(\key_mem[12][15] ), .IN2(n6633), .IN3(\key_mem[13][15] ), .IN4(
          n6618), .IN5(n5666), .Q(n5669));
   AO22X1 U6323 (.IN1(\key_mem[7][15] ), .IN2(n6663), .IN3(\key_mem[2][15] ), .IN4(n6648)
          , .Q(n5667));
   AO221X1 U6324 (.IN1(\key_mem[0][15] ), .IN2(n6693), .IN3(\key_mem[1][15] ), .IN4(n6678)
          , .IN5(n5667), .Q(n5668));
   OR4X1 U6325 (.IN1(n5671), .IN2(n5670), .IN3(n5669), .IN4(n5668), .Q(round_key[15]));
   AO22X1 U6326 (.IN1(\key_mem[11][16] ), .IN2(n6498), .IN3(\key_mem[6][16] ), .IN4(n6483)
          , .Q(n5672));
   AO221X1 U6327 (.IN1(\key_mem[4][16] ), .IN2(n6528), .IN3(\key_mem[5][16] ), .IN4(n6513)
          , .IN5(n5672), .Q(n5678));
   AO222X1 U6328 (.IN1(\key_mem[9][16] ), .IN2(n6573), .IN3(\key_mem[8][16] ), .IN4(n6558)
          , .IN5(\key_mem[10][16] ), .IN6(n6543), .Q(n5677));
   AO22X1 U6329 (.IN1(\key_mem[3][16] ), .IN2(n6603), .IN3(\key_mem[14][16] ), .IN4(n6588)
          , .Q(n5673));
   AO221X1 U6330 (.IN1(\key_mem[12][16] ), .IN2(n6633), .IN3(\key_mem[13][16] ), .IN4(
          n6618), .IN5(n5673), .Q(n5676));
   AO22X1 U6331 (.IN1(\key_mem[7][16] ), .IN2(n6663), .IN3(\key_mem[2][16] ), .IN4(n6648)
          , .Q(n5674));
   AO221X1 U6332 (.IN1(\key_mem[0][16] ), .IN2(n6693), .IN3(\key_mem[1][16] ), .IN4(n6678)
          , .IN5(n5674), .Q(n5675));
   OR4X1 U6333 (.IN1(n5678), .IN2(n5677), .IN3(n5676), .IN4(n5675), .Q(round_key[16]));
   AO22X1 U6334 (.IN1(\key_mem[11][17] ), .IN2(n6498), .IN3(\key_mem[6][17] ), .IN4(n6483)
          , .Q(n5679));
   AO221X1 U6335 (.IN1(\key_mem[4][17] ), .IN2(n6528), .IN3(\key_mem[5][17] ), .IN4(n6513)
          , .IN5(n5679), .Q(n5685));
   AO222X1 U6336 (.IN1(\key_mem[9][17] ), .IN2(n6573), .IN3(\key_mem[8][17] ), .IN4(n6558)
          , .IN5(\key_mem[10][17] ), .IN6(n6543), .Q(n5684));
   AO22X1 U6337 (.IN1(\key_mem[3][17] ), .IN2(n6603), .IN3(\key_mem[14][17] ), .IN4(n6588)
          , .Q(n5680));
   AO221X1 U6338 (.IN1(\key_mem[12][17] ), .IN2(n6633), .IN3(\key_mem[13][17] ), .IN4(
          n6618), .IN5(n5680), .Q(n5683));
   AO22X1 U6339 (.IN1(\key_mem[7][17] ), .IN2(n6663), .IN3(\key_mem[2][17] ), .IN4(n6648)
          , .Q(n5681));
   AO221X1 U6340 (.IN1(\key_mem[0][17] ), .IN2(n6693), .IN3(\key_mem[1][17] ), .IN4(n6678)
          , .IN5(n5681), .Q(n5682));
   OR4X1 U6341 (.IN1(n5685), .IN2(n5684), .IN3(n5683), .IN4(n5682), .Q(round_key[17]));
   AO22X1 U6342 (.IN1(\key_mem[11][18] ), .IN2(n6498), .IN3(\key_mem[6][18] ), .IN4(n6483)
          , .Q(n5686));
   AO221X1 U6343 (.IN1(\key_mem[4][18] ), .IN2(n6528), .IN3(\key_mem[5][18] ), .IN4(n6513)
          , .IN5(n5686), .Q(n5692));
   AO222X1 U6344 (.IN1(\key_mem[9][18] ), .IN2(n6573), .IN3(\key_mem[8][18] ), .IN4(n6558)
          , .IN5(\key_mem[10][18] ), .IN6(n6543), .Q(n5691));
   AO22X1 U6345 (.IN1(\key_mem[3][18] ), .IN2(n6603), .IN3(\key_mem[14][18] ), .IN4(n6588)
          , .Q(n5687));
   AO221X1 U6346 (.IN1(\key_mem[12][18] ), .IN2(n6633), .IN3(\key_mem[13][18] ), .IN4(
          n6618), .IN5(n5687), .Q(n5690));
   AO22X1 U6347 (.IN1(\key_mem[7][18] ), .IN2(n6663), .IN3(\key_mem[2][18] ), .IN4(n6648)
          , .Q(n5688));
   AO221X1 U6348 (.IN1(\key_mem[0][18] ), .IN2(n6693), .IN3(\key_mem[1][18] ), .IN4(n6678)
          , .IN5(n5688), .Q(n5689));
   OR4X1 U6349 (.IN1(n5692), .IN2(n5691), .IN3(n5690), .IN4(n5689), .Q(round_key[18]));
   AO22X1 U6350 (.IN1(\key_mem[11][19] ), .IN2(n6498), .IN3(\key_mem[6][19] ), .IN4(n6483)
          , .Q(n5693));
   AO221X1 U6351 (.IN1(\key_mem[4][19] ), .IN2(n6528), .IN3(\key_mem[5][19] ), .IN4(n6513)
          , .IN5(n5693), .Q(n5699));
   AO222X1 U6352 (.IN1(\key_mem[9][19] ), .IN2(n6573), .IN3(\key_mem[8][19] ), .IN4(n6558)
          , .IN5(\key_mem[10][19] ), .IN6(n6543), .Q(n5698));
   AO22X1 U6353 (.IN1(\key_mem[3][19] ), .IN2(n6603), .IN3(\key_mem[14][19] ), .IN4(n6588)
          , .Q(n5694));
   AO221X1 U6354 (.IN1(\key_mem[12][19] ), .IN2(n6633), .IN3(\key_mem[13][19] ), .IN4(
          n6618), .IN5(n5694), .Q(n5697));
   AO22X1 U6355 (.IN1(\key_mem[7][19] ), .IN2(n6663), .IN3(\key_mem[2][19] ), .IN4(n6648)
          , .Q(n5695));
   AO221X1 U6356 (.IN1(\key_mem[0][19] ), .IN2(n6693), .IN3(\key_mem[1][19] ), .IN4(n6678)
          , .IN5(n5695), .Q(n5696));
   OR4X1 U6357 (.IN1(n5699), .IN2(n5698), .IN3(n5697), .IN4(n5696), .Q(round_key[19]));
   AO22X1 U6358 (.IN1(\key_mem[11][20] ), .IN2(n6498), .IN3(\key_mem[6][20] ), .IN4(n6483)
          , .Q(n5700));
   AO221X1 U6359 (.IN1(\key_mem[4][20] ), .IN2(n6528), .IN3(\key_mem[5][20] ), .IN4(n6513)
          , .IN5(n5700), .Q(n5706));
   AO222X1 U6360 (.IN1(\key_mem[9][20] ), .IN2(n6573), .IN3(\key_mem[8][20] ), .IN4(n6558)
          , .IN5(\key_mem[10][20] ), .IN6(n6543), .Q(n5705));
   AO22X1 U6361 (.IN1(\key_mem[3][20] ), .IN2(n6603), .IN3(\key_mem[14][20] ), .IN4(n6588)
          , .Q(n5701));
   AO221X1 U6362 (.IN1(\key_mem[12][20] ), .IN2(n6633), .IN3(\key_mem[13][20] ), .IN4(
          n6618), .IN5(n5701), .Q(n5704));
   AO22X1 U6363 (.IN1(\key_mem[7][20] ), .IN2(n6663), .IN3(\key_mem[2][20] ), .IN4(n6648)
          , .Q(n5702));
   AO221X1 U6364 (.IN1(\key_mem[0][20] ), .IN2(n6693), .IN3(\key_mem[1][20] ), .IN4(n6678)
          , .IN5(n5702), .Q(n5703));
   OR4X1 U6365 (.IN1(n5706), .IN2(n5705), .IN3(n5704), .IN4(n5703), .Q(round_key[20]));
   AO22X1 U6366 (.IN1(\key_mem[11][21] ), .IN2(n6498), .IN3(\key_mem[6][21] ), .IN4(n6483)
          , .Q(n5707));
   AO221X1 U6367 (.IN1(\key_mem[4][21] ), .IN2(n6528), .IN3(\key_mem[5][21] ), .IN4(n6513)
          , .IN5(n5707), .Q(n5713));
   AO222X1 U6368 (.IN1(\key_mem[9][21] ), .IN2(n6573), .IN3(\key_mem[8][21] ), .IN4(n6558)
          , .IN5(\key_mem[10][21] ), .IN6(n6543), .Q(n5712));
   AO22X1 U6369 (.IN1(\key_mem[3][21] ), .IN2(n6603), .IN3(\key_mem[14][21] ), .IN4(n6588)
          , .Q(n5708));
   AO221X1 U6370 (.IN1(\key_mem[12][21] ), .IN2(n6633), .IN3(\key_mem[13][21] ), .IN4(
          n6618), .IN5(n5708), .Q(n5711));
   AO22X1 U6371 (.IN1(\key_mem[7][21] ), .IN2(n6663), .IN3(\key_mem[2][21] ), .IN4(n6648)
          , .Q(n5709));
   AO221X1 U6372 (.IN1(\key_mem[0][21] ), .IN2(n6693), .IN3(\key_mem[1][21] ), .IN4(n6678)
          , .IN5(n5709), .Q(n5710));
   OR4X1 U6373 (.IN1(n5713), .IN2(n5712), .IN3(n5711), .IN4(n5710), .Q(round_key[21]));
   AO22X1 U6374 (.IN1(\key_mem[11][22] ), .IN2(n6498), .IN3(\key_mem[6][22] ), .IN4(n6483)
          , .Q(n5714));
   AO221X1 U6375 (.IN1(\key_mem[4][22] ), .IN2(n6528), .IN3(\key_mem[5][22] ), .IN4(n6513)
          , .IN5(n5714), .Q(n5720));
   AO222X1 U6376 (.IN1(\key_mem[9][22] ), .IN2(n6573), .IN3(\key_mem[8][22] ), .IN4(n6558)
          , .IN5(\key_mem[10][22] ), .IN6(n6543), .Q(n5719));
   AO22X1 U6377 (.IN1(\key_mem[3][22] ), .IN2(n6603), .IN3(\key_mem[14][22] ), .IN4(n6588)
          , .Q(n5715));
   AO221X1 U6378 (.IN1(\key_mem[12][22] ), .IN2(n6633), .IN3(\key_mem[13][22] ), .IN4(
          n6618), .IN5(n5715), .Q(n5718));
   AO22X1 U6379 (.IN1(\key_mem[7][22] ), .IN2(n6663), .IN3(\key_mem[2][22] ), .IN4(n6648)
          , .Q(n5716));
   AO221X1 U6380 (.IN1(\key_mem[0][22] ), .IN2(n6693), .IN3(\key_mem[1][22] ), .IN4(n6678)
          , .IN5(n5716), .Q(n5717));
   OR4X1 U6381 (.IN1(n5720), .IN2(n5719), .IN3(n5718), .IN4(n5717), .Q(round_key[22]));
   AO22X1 U6382 (.IN1(\key_mem[11][23] ), .IN2(n6498), .IN3(\key_mem[6][23] ), .IN4(n6483)
          , .Q(n5721));
   AO221X1 U6383 (.IN1(\key_mem[4][23] ), .IN2(n6528), .IN3(\key_mem[5][23] ), .IN4(n6513)
          , .IN5(n5721), .Q(n5727));
   AO222X1 U6384 (.IN1(\key_mem[9][23] ), .IN2(n6573), .IN3(\key_mem[8][23] ), .IN4(n6558)
          , .IN5(\key_mem[10][23] ), .IN6(n6543), .Q(n5726));
   AO22X1 U6385 (.IN1(\key_mem[3][23] ), .IN2(n6603), .IN3(\key_mem[14][23] ), .IN4(n6588)
          , .Q(n5722));
   AO221X1 U6386 (.IN1(\key_mem[12][23] ), .IN2(n6633), .IN3(\key_mem[13][23] ), .IN4(
          n6618), .IN5(n5722), .Q(n5725));
   AO22X1 U6387 (.IN1(\key_mem[7][23] ), .IN2(n6663), .IN3(\key_mem[2][23] ), .IN4(n6648)
          , .Q(n5723));
   AO221X1 U6388 (.IN1(\key_mem[0][23] ), .IN2(n6693), .IN3(\key_mem[1][23] ), .IN4(n6678)
          , .IN5(n5723), .Q(n5724));
   OR4X1 U6389 (.IN1(n5727), .IN2(n5726), .IN3(n5725), .IN4(n5724), .Q(round_key[23]));
   AO22X1 U6390 (.IN1(\key_mem[11][24] ), .IN2(n6497), .IN3(\key_mem[6][24] ), .IN4(n6482)
          , .Q(n5728));
   AO221X1 U6391 (.IN1(\key_mem[4][24] ), .IN2(n6527), .IN3(\key_mem[5][24] ), .IN4(n6512)
          , .IN5(n5728), .Q(n5734));
   AO222X1 U6392 (.IN1(\key_mem[9][24] ), .IN2(n6572), .IN3(\key_mem[8][24] ), .IN4(n6557)
          , .IN5(\key_mem[10][24] ), .IN6(n6542), .Q(n5733));
   AO22X1 U6393 (.IN1(\key_mem[3][24] ), .IN2(n6602), .IN3(\key_mem[14][24] ), .IN4(n6587)
          , .Q(n5729));
   AO221X1 U6394 (.IN1(\key_mem[12][24] ), .IN2(n6632), .IN3(\key_mem[13][24] ), .IN4(
          n6617), .IN5(n5729), .Q(n5732));
   AO22X1 U6395 (.IN1(\key_mem[7][24] ), .IN2(n6662), .IN3(\key_mem[2][24] ), .IN4(n6647)
          , .Q(n5730));
   AO221X1 U6396 (.IN1(\key_mem[0][24] ), .IN2(n6692), .IN3(\key_mem[1][24] ), .IN4(n6677)
          , .IN5(n5730), .Q(n5731));
   OR4X1 U6397 (.IN1(n5734), .IN2(n5733), .IN3(n5732), .IN4(n5731), .Q(round_key[24]));
   AO22X1 U6398 (.IN1(\key_mem[11][25] ), .IN2(n6497), .IN3(\key_mem[6][25] ), .IN4(n6482)
          , .Q(n5735));
   AO221X1 U6399 (.IN1(\key_mem[4][25] ), .IN2(n6527), .IN3(\key_mem[5][25] ), .IN4(n6512)
          , .IN5(n5735), .Q(n5741));
   AO222X1 U6400 (.IN1(\key_mem[9][25] ), .IN2(n6572), .IN3(\key_mem[8][25] ), .IN4(n6557)
          , .IN5(\key_mem[10][25] ), .IN6(n6542), .Q(n5740));
   AO22X1 U6401 (.IN1(\key_mem[3][25] ), .IN2(n6602), .IN3(\key_mem[14][25] ), .IN4(n6587)
          , .Q(n5736));
   AO221X1 U6402 (.IN1(\key_mem[12][25] ), .IN2(n6632), .IN3(\key_mem[13][25] ), .IN4(
          n6617), .IN5(n5736), .Q(n5739));
   AO22X1 U6403 (.IN1(\key_mem[7][25] ), .IN2(n6662), .IN3(\key_mem[2][25] ), .IN4(n6647)
          , .Q(n5737));
   AO221X1 U6404 (.IN1(\key_mem[0][25] ), .IN2(n6692), .IN3(\key_mem[1][25] ), .IN4(n6677)
          , .IN5(n5737), .Q(n5738));
   OR4X1 U6405 (.IN1(n5741), .IN2(n5740), .IN3(n5739), .IN4(n5738), .Q(round_key[25]));
   AO22X1 U6406 (.IN1(\key_mem[11][26] ), .IN2(n6497), .IN3(\key_mem[6][26] ), .IN4(n6482)
          , .Q(n5742));
   AO221X1 U6407 (.IN1(\key_mem[4][26] ), .IN2(n6527), .IN3(\key_mem[5][26] ), .IN4(n6512)
          , .IN5(n5742), .Q(n5748));
   AO222X1 U6408 (.IN1(\key_mem[9][26] ), .IN2(n6572), .IN3(\key_mem[8][26] ), .IN4(n6557)
          , .IN5(\key_mem[10][26] ), .IN6(n6542), .Q(n5747));
   AO22X1 U6409 (.IN1(\key_mem[3][26] ), .IN2(n6602), .IN3(\key_mem[14][26] ), .IN4(n6587)
          , .Q(n5743));
   AO221X1 U6410 (.IN1(\key_mem[12][26] ), .IN2(n6632), .IN3(\key_mem[13][26] ), .IN4(
          n6617), .IN5(n5743), .Q(n5746));
   AO22X1 U6411 (.IN1(\key_mem[7][26] ), .IN2(n6662), .IN3(\key_mem[2][26] ), .IN4(n6647)
          , .Q(n5744));
   AO221X1 U6412 (.IN1(\key_mem[0][26] ), .IN2(n6692), .IN3(\key_mem[1][26] ), .IN4(n6677)
          , .IN5(n5744), .Q(n5745));
   OR4X1 U6413 (.IN1(n5748), .IN2(n5747), .IN3(n5746), .IN4(n5745), .Q(round_key[26]));
   AO22X1 U6414 (.IN1(\key_mem[11][27] ), .IN2(n6497), .IN3(\key_mem[6][27] ), .IN4(n6482)
          , .Q(n5749));
   AO221X1 U6415 (.IN1(\key_mem[4][27] ), .IN2(n6527), .IN3(\key_mem[5][27] ), .IN4(n6512)
          , .IN5(n5749), .Q(n5755));
   AO222X1 U6416 (.IN1(\key_mem[9][27] ), .IN2(n6572), .IN3(\key_mem[8][27] ), .IN4(n6557)
          , .IN5(\key_mem[10][27] ), .IN6(n6542), .Q(n5754));
   AO22X1 U6417 (.IN1(\key_mem[3][27] ), .IN2(n6602), .IN3(\key_mem[14][27] ), .IN4(n6587)
          , .Q(n5750));
   AO221X1 U6418 (.IN1(\key_mem[12][27] ), .IN2(n6632), .IN3(\key_mem[13][27] ), .IN4(
          n6617), .IN5(n5750), .Q(n5753));
   AO22X1 U6419 (.IN1(\key_mem[7][27] ), .IN2(n6662), .IN3(\key_mem[2][27] ), .IN4(n6647)
          , .Q(n5751));
   AO221X1 U6420 (.IN1(\key_mem[0][27] ), .IN2(n6692), .IN3(\key_mem[1][27] ), .IN4(n6677)
          , .IN5(n5751), .Q(n5752));
   OR4X1 U6421 (.IN1(n5755), .IN2(n5754), .IN3(n5753), .IN4(n5752), .Q(round_key[27]));
   AO22X1 U6422 (.IN1(\key_mem[11][28] ), .IN2(n6497), .IN3(\key_mem[6][28] ), .IN4(n6482)
          , .Q(n5756));
   AO221X1 U6423 (.IN1(\key_mem[4][28] ), .IN2(n6527), .IN3(\key_mem[5][28] ), .IN4(n6512)
          , .IN5(n5756), .Q(n5762));
   AO222X1 U6424 (.IN1(\key_mem[9][28] ), .IN2(n6572), .IN3(\key_mem[8][28] ), .IN4(n6557)
          , .IN5(\key_mem[10][28] ), .IN6(n6542), .Q(n5761));
   AO22X1 U6425 (.IN1(\key_mem[3][28] ), .IN2(n6602), .IN3(\key_mem[14][28] ), .IN4(n6587)
          , .Q(n5757));
   AO221X1 U6426 (.IN1(\key_mem[12][28] ), .IN2(n6632), .IN3(\key_mem[13][28] ), .IN4(
          n6617), .IN5(n5757), .Q(n5760));
   AO22X1 U6427 (.IN1(\key_mem[7][28] ), .IN2(n6662), .IN3(\key_mem[2][28] ), .IN4(n6647)
          , .Q(n5758));
   AO221X1 U6428 (.IN1(\key_mem[0][28] ), .IN2(n6692), .IN3(\key_mem[1][28] ), .IN4(n6677)
          , .IN5(n5758), .Q(n5759));
   OR4X1 U6429 (.IN1(n5762), .IN2(n5761), .IN3(n5760), .IN4(n5759), .Q(round_key[28]));
   AO22X1 U6430 (.IN1(\key_mem[11][29] ), .IN2(n6497), .IN3(\key_mem[6][29] ), .IN4(n6482)
          , .Q(n5763));
   AO221X1 U6431 (.IN1(\key_mem[4][29] ), .IN2(n6527), .IN3(\key_mem[5][29] ), .IN4(n6512)
          , .IN5(n5763), .Q(n5769));
   AO222X1 U6432 (.IN1(\key_mem[9][29] ), .IN2(n6572), .IN3(\key_mem[8][29] ), .IN4(n6557)
          , .IN5(\key_mem[10][29] ), .IN6(n6542), .Q(n5768));
   AO22X1 U6433 (.IN1(\key_mem[3][29] ), .IN2(n6602), .IN3(\key_mem[14][29] ), .IN4(n6587)
          , .Q(n5764));
   AO221X1 U6434 (.IN1(\key_mem[12][29] ), .IN2(n6632), .IN3(\key_mem[13][29] ), .IN4(
          n6617), .IN5(n5764), .Q(n5767));
   AO22X1 U6435 (.IN1(\key_mem[7][29] ), .IN2(n6662), .IN3(\key_mem[2][29] ), .IN4(n6647)
          , .Q(n5765));
   AO221X1 U6436 (.IN1(\key_mem[0][29] ), .IN2(n6692), .IN3(\key_mem[1][29] ), .IN4(n6677)
          , .IN5(n5765), .Q(n5766));
   OR4X1 U6437 (.IN1(n5769), .IN2(n5768), .IN3(n5767), .IN4(n5766), .Q(round_key[29]));
   AO22X1 U6438 (.IN1(\key_mem[11][30] ), .IN2(n6497), .IN3(\key_mem[6][30] ), .IN4(n6482)
          , .Q(n5770));
   AO221X1 U6439 (.IN1(\key_mem[4][30] ), .IN2(n6527), .IN3(\key_mem[5][30] ), .IN4(n6512)
          , .IN5(n5770), .Q(n5776));
   AO222X1 U6440 (.IN1(\key_mem[9][30] ), .IN2(n6572), .IN3(\key_mem[8][30] ), .IN4(n6557)
          , .IN5(\key_mem[10][30] ), .IN6(n6542), .Q(n5775));
   AO22X1 U6441 (.IN1(\key_mem[3][30] ), .IN2(n6602), .IN3(\key_mem[14][30] ), .IN4(n6587)
          , .Q(n5771));
   AO221X1 U6442 (.IN1(\key_mem[12][30] ), .IN2(n6632), .IN3(\key_mem[13][30] ), .IN4(
          n6617), .IN5(n5771), .Q(n5774));
   AO22X1 U6443 (.IN1(\key_mem[7][30] ), .IN2(n6662), .IN3(\key_mem[2][30] ), .IN4(n6647)
          , .Q(n5772));
   AO221X1 U6444 (.IN1(\key_mem[0][30] ), .IN2(n6692), .IN3(\key_mem[1][30] ), .IN4(n6677)
          , .IN5(n5772), .Q(n5773));
   OR4X1 U6445 (.IN1(n5776), .IN2(n5775), .IN3(n5774), .IN4(n5773), .Q(round_key[30]));
   AO22X1 U6446 (.IN1(\key_mem[11][31] ), .IN2(n6497), .IN3(\key_mem[6][31] ), .IN4(n6482)
          , .Q(n5777));
   AO221X1 U6447 (.IN1(\key_mem[4][31] ), .IN2(n6527), .IN3(\key_mem[5][31] ), .IN4(n6512)
          , .IN5(n5777), .Q(n5783));
   AO222X1 U6448 (.IN1(\key_mem[9][31] ), .IN2(n6572), .IN3(\key_mem[8][31] ), .IN4(n6557)
          , .IN5(\key_mem[10][31] ), .IN6(n6542), .Q(n5782));
   AO22X1 U6449 (.IN1(\key_mem[3][31] ), .IN2(n6602), .IN3(\key_mem[14][31] ), .IN4(n6587)
          , .Q(n5778));
   AO221X1 U6450 (.IN1(\key_mem[12][31] ), .IN2(n6632), .IN3(\key_mem[13][31] ), .IN4(
          n6617), .IN5(n5778), .Q(n5781));
   AO22X1 U6451 (.IN1(\key_mem[7][31] ), .IN2(n6662), .IN3(\key_mem[2][31] ), .IN4(n6647)
          , .Q(n5779));
   AO221X1 U6452 (.IN1(\key_mem[0][31] ), .IN2(n6692), .IN3(\key_mem[1][31] ), .IN4(n6677)
          , .IN5(n5779), .Q(n5780));
   OR4X1 U6453 (.IN1(n5783), .IN2(n5782), .IN3(n5781), .IN4(n5780), .Q(round_key[31]));
   AO22X1 U6454 (.IN1(\key_mem[11][32] ), .IN2(n6497), .IN3(\key_mem[6][32] ), .IN4(n6482)
          , .Q(n5784));
   AO221X1 U6455 (.IN1(\key_mem[4][32] ), .IN2(n6527), .IN3(\key_mem[5][32] ), .IN4(n6512)
          , .IN5(n5784), .Q(n5790));
   AO222X1 U6456 (.IN1(\key_mem[9][32] ), .IN2(n6572), .IN3(\key_mem[8][32] ), .IN4(n6557)
          , .IN5(\key_mem[10][32] ), .IN6(n6542), .Q(n5789));
   AO22X1 U6457 (.IN1(\key_mem[3][32] ), .IN2(n6602), .IN3(\key_mem[14][32] ), .IN4(n6587)
          , .Q(n5785));
   AO221X1 U6458 (.IN1(\key_mem[12][32] ), .IN2(n6632), .IN3(\key_mem[13][32] ), .IN4(
          n6617), .IN5(n5785), .Q(n5788));
   AO22X1 U6459 (.IN1(\key_mem[7][32] ), .IN2(n6662), .IN3(\key_mem[2][32] ), .IN4(n6647)
          , .Q(n5786));
   AO221X1 U6460 (.IN1(\key_mem[0][32] ), .IN2(n6692), .IN3(\key_mem[1][32] ), .IN4(n6677)
          , .IN5(n5786), .Q(n5787));
   OR4X1 U6461 (.IN1(n5790), .IN2(n5789), .IN3(n5788), .IN4(n5787), .Q(round_key[32]));
   AO22X1 U6462 (.IN1(\key_mem[11][33] ), .IN2(n6497), .IN3(\key_mem[6][33] ), .IN4(n6482)
          , .Q(n5791));
   AO221X1 U6463 (.IN1(\key_mem[4][33] ), .IN2(n6527), .IN3(\key_mem[5][33] ), .IN4(n6512)
          , .IN5(n5791), .Q(n5797));
   AO222X1 U6464 (.IN1(\key_mem[9][33] ), .IN2(n6572), .IN3(\key_mem[8][33] ), .IN4(n6557)
          , .IN5(\key_mem[10][33] ), .IN6(n6542), .Q(n5796));
   AO22X1 U6465 (.IN1(\key_mem[3][33] ), .IN2(n6602), .IN3(\key_mem[14][33] ), .IN4(n6587)
          , .Q(n5792));
   AO221X1 U6466 (.IN1(\key_mem[12][33] ), .IN2(n6632), .IN3(\key_mem[13][33] ), .IN4(
          n6617), .IN5(n5792), .Q(n5795));
   AO22X1 U6467 (.IN1(\key_mem[7][33] ), .IN2(n6662), .IN3(\key_mem[2][33] ), .IN4(n6647)
          , .Q(n5793));
   AO221X1 U6468 (.IN1(\key_mem[0][33] ), .IN2(n6692), .IN3(\key_mem[1][33] ), .IN4(n6677)
          , .IN5(n5793), .Q(n5794));
   OR4X1 U6469 (.IN1(n5797), .IN2(n5796), .IN3(n5795), .IN4(n5794), .Q(round_key[33]));
   AO22X1 U6470 (.IN1(\key_mem[11][34] ), .IN2(n6497), .IN3(\key_mem[6][34] ), .IN4(n6482)
          , .Q(n5798));
   AO221X1 U6471 (.IN1(\key_mem[4][34] ), .IN2(n6527), .IN3(\key_mem[5][34] ), .IN4(n6512)
          , .IN5(n5798), .Q(n5804));
   AO222X1 U6472 (.IN1(\key_mem[9][34] ), .IN2(n6572), .IN3(\key_mem[8][34] ), .IN4(n6557)
          , .IN5(\key_mem[10][34] ), .IN6(n6542), .Q(n5803));
   AO22X1 U6473 (.IN1(\key_mem[3][34] ), .IN2(n6602), .IN3(\key_mem[14][34] ), .IN4(n6587)
          , .Q(n5799));
   AO221X1 U6474 (.IN1(\key_mem[12][34] ), .IN2(n6632), .IN3(\key_mem[13][34] ), .IN4(
          n6617), .IN5(n5799), .Q(n5802));
   AO22X1 U6475 (.IN1(\key_mem[7][34] ), .IN2(n6662), .IN3(\key_mem[2][34] ), .IN4(n6647)
          , .Q(n5800));
   AO221X1 U6476 (.IN1(\key_mem[0][34] ), .IN2(n6692), .IN3(\key_mem[1][34] ), .IN4(n6677)
          , .IN5(n5800), .Q(n5801));
   OR4X1 U6477 (.IN1(n5804), .IN2(n5803), .IN3(n5802), .IN4(n5801), .Q(round_key[34]));
   AO22X1 U6478 (.IN1(\key_mem[11][35] ), .IN2(n6497), .IN3(\key_mem[6][35] ), .IN4(n6482)
          , .Q(n5805));
   AO221X1 U6479 (.IN1(\key_mem[4][35] ), .IN2(n6527), .IN3(\key_mem[5][35] ), .IN4(n6512)
          , .IN5(n5805), .Q(n5811));
   AO222X1 U6480 (.IN1(\key_mem[9][35] ), .IN2(n6572), .IN3(\key_mem[8][35] ), .IN4(n6557)
          , .IN5(\key_mem[10][35] ), .IN6(n6542), .Q(n5810));
   AO22X1 U6481 (.IN1(\key_mem[3][35] ), .IN2(n6602), .IN3(\key_mem[14][35] ), .IN4(n6587)
          , .Q(n5806));
   AO221X1 U6482 (.IN1(\key_mem[12][35] ), .IN2(n6632), .IN3(\key_mem[13][35] ), .IN4(
          n6617), .IN5(n5806), .Q(n5809));
   AO22X1 U6483 (.IN1(\key_mem[7][35] ), .IN2(n6662), .IN3(\key_mem[2][35] ), .IN4(n6647)
          , .Q(n5807));
   AO221X1 U6484 (.IN1(\key_mem[0][35] ), .IN2(n6692), .IN3(\key_mem[1][35] ), .IN4(n6677)
          , .IN5(n5807), .Q(n5808));
   OR4X1 U6485 (.IN1(n5811), .IN2(n5810), .IN3(n5809), .IN4(n5808), .Q(round_key[35]));
   AO22X1 U6486 (.IN1(\key_mem[11][36] ), .IN2(n6496), .IN3(\key_mem[6][36] ), .IN4(n6481)
          , .Q(n5812));
   AO221X1 U6487 (.IN1(\key_mem[4][36] ), .IN2(n6526), .IN3(\key_mem[5][36] ), .IN4(n6511)
          , .IN5(n5812), .Q(n5818));
   AO222X1 U6488 (.IN1(\key_mem[9][36] ), .IN2(n6571), .IN3(\key_mem[8][36] ), .IN4(n6556)
          , .IN5(\key_mem[10][36] ), .IN6(n6541), .Q(n5817));
   AO22X1 U6489 (.IN1(\key_mem[3][36] ), .IN2(n6601), .IN3(\key_mem[14][36] ), .IN4(n6586)
          , .Q(n5813));
   AO221X1 U6490 (.IN1(\key_mem[12][36] ), .IN2(n6631), .IN3(\key_mem[13][36] ), .IN4(
          n6616), .IN5(n5813), .Q(n5816));
   AO22X1 U6491 (.IN1(\key_mem[7][36] ), .IN2(n6661), .IN3(\key_mem[2][36] ), .IN4(n6646)
          , .Q(n5814));
   AO221X1 U6492 (.IN1(\key_mem[0][36] ), .IN2(n6691), .IN3(\key_mem[1][36] ), .IN4(n6676)
          , .IN5(n5814), .Q(n5815));
   OR4X1 U6493 (.IN1(n5818), .IN2(n5817), .IN3(n5816), .IN4(n5815), .Q(round_key[36]));
   AO22X1 U6494 (.IN1(\key_mem[11][37] ), .IN2(n6496), .IN3(\key_mem[6][37] ), .IN4(n6481)
          , .Q(n5819));
   AO221X1 U6495 (.IN1(\key_mem[4][37] ), .IN2(n6526), .IN3(\key_mem[5][37] ), .IN4(n6511)
          , .IN5(n5819), .Q(n5825));
   AO222X1 U6496 (.IN1(\key_mem[9][37] ), .IN2(n6571), .IN3(\key_mem[8][37] ), .IN4(n6556)
          , .IN5(\key_mem[10][37] ), .IN6(n6541), .Q(n5824));
   AO22X1 U6497 (.IN1(\key_mem[3][37] ), .IN2(n6601), .IN3(\key_mem[14][37] ), .IN4(n6586)
          , .Q(n5820));
   AO221X1 U6498 (.IN1(\key_mem[12][37] ), .IN2(n6631), .IN3(\key_mem[13][37] ), .IN4(
          n6616), .IN5(n5820), .Q(n5823));
   AO22X1 U6499 (.IN1(\key_mem[7][37] ), .IN2(n6661), .IN3(\key_mem[2][37] ), .IN4(n6646)
          , .Q(n5821));
   AO221X1 U6500 (.IN1(\key_mem[0][37] ), .IN2(n6691), .IN3(\key_mem[1][37] ), .IN4(n6676)
          , .IN5(n5821), .Q(n5822));
   OR4X1 U6501 (.IN1(n5825), .IN2(n5824), .IN3(n5823), .IN4(n5822), .Q(round_key[37]));
   AO22X1 U6502 (.IN1(\key_mem[11][38] ), .IN2(n6496), .IN3(\key_mem[6][38] ), .IN4(n6481)
          , .Q(n5826));
   AO221X1 U6503 (.IN1(\key_mem[4][38] ), .IN2(n6526), .IN3(\key_mem[5][38] ), .IN4(n6511)
          , .IN5(n5826), .Q(n5832));
   AO222X1 U6504 (.IN1(\key_mem[9][38] ), .IN2(n6571), .IN3(\key_mem[8][38] ), .IN4(n6556)
          , .IN5(\key_mem[10][38] ), .IN6(n6541), .Q(n5831));
   AO22X1 U6505 (.IN1(\key_mem[3][38] ), .IN2(n6601), .IN3(\key_mem[14][38] ), .IN4(n6586)
          , .Q(n5827));
   AO221X1 U6506 (.IN1(\key_mem[12][38] ), .IN2(n6631), .IN3(\key_mem[13][38] ), .IN4(
          n6616), .IN5(n5827), .Q(n5830));
   AO22X1 U6507 (.IN1(\key_mem[7][38] ), .IN2(n6661), .IN3(\key_mem[2][38] ), .IN4(n6646)
          , .Q(n5828));
   AO221X1 U6508 (.IN1(\key_mem[0][38] ), .IN2(n6691), .IN3(\key_mem[1][38] ), .IN4(n6676)
          , .IN5(n5828), .Q(n5829));
   OR4X1 U6509 (.IN1(n5832), .IN2(n5831), .IN3(n5830), .IN4(n5829), .Q(round_key[38]));
   AO22X1 U6510 (.IN1(\key_mem[11][39] ), .IN2(n6496), .IN3(\key_mem[6][39] ), .IN4(n6481)
          , .Q(n5833));
   AO221X1 U6511 (.IN1(\key_mem[4][39] ), .IN2(n6526), .IN3(\key_mem[5][39] ), .IN4(n6511)
          , .IN5(n5833), .Q(n5839));
   AO222X1 U6512 (.IN1(\key_mem[9][39] ), .IN2(n6571), .IN3(\key_mem[8][39] ), .IN4(n6556)
          , .IN5(\key_mem[10][39] ), .IN6(n6541), .Q(n5838));
   AO22X1 U6513 (.IN1(\key_mem[3][39] ), .IN2(n6601), .IN3(\key_mem[14][39] ), .IN4(n6586)
          , .Q(n5834));
   AO221X1 U6514 (.IN1(\key_mem[12][39] ), .IN2(n6631), .IN3(\key_mem[13][39] ), .IN4(
          n6616), .IN5(n5834), .Q(n5837));
   AO22X1 U6515 (.IN1(\key_mem[7][39] ), .IN2(n6661), .IN3(\key_mem[2][39] ), .IN4(n6646)
          , .Q(n5835));
   AO221X1 U6516 (.IN1(\key_mem[0][39] ), .IN2(n6691), .IN3(\key_mem[1][39] ), .IN4(n6676)
          , .IN5(n5835), .Q(n5836));
   OR4X1 U6517 (.IN1(n5839), .IN2(n5838), .IN3(n5837), .IN4(n5836), .Q(round_key[39]));
   AO22X1 U6518 (.IN1(\key_mem[11][40] ), .IN2(n6496), .IN3(\key_mem[6][40] ), .IN4(n6481)
          , .Q(n5840));
   AO221X1 U6519 (.IN1(\key_mem[4][40] ), .IN2(n6526), .IN3(\key_mem[5][40] ), .IN4(n6511)
          , .IN5(n5840), .Q(n5846));
   AO222X1 U6520 (.IN1(\key_mem[9][40] ), .IN2(n6571), .IN3(\key_mem[8][40] ), .IN4(n6556)
          , .IN5(\key_mem[10][40] ), .IN6(n6541), .Q(n5845));
   AO22X1 U6521 (.IN1(\key_mem[3][40] ), .IN2(n6601), .IN3(\key_mem[14][40] ), .IN4(n6586)
          , .Q(n5841));
   AO221X1 U6522 (.IN1(\key_mem[12][40] ), .IN2(n6631), .IN3(\key_mem[13][40] ), .IN4(
          n6616), .IN5(n5841), .Q(n5844));
   AO22X1 U6523 (.IN1(\key_mem[7][40] ), .IN2(n6661), .IN3(\key_mem[2][40] ), .IN4(n6646)
          , .Q(n5842));
   AO221X1 U6524 (.IN1(\key_mem[0][40] ), .IN2(n6691), .IN3(\key_mem[1][40] ), .IN4(n6676)
          , .IN5(n5842), .Q(n5843));
   OR4X1 U6525 (.IN1(n5846), .IN2(n5845), .IN3(n5844), .IN4(n5843), .Q(round_key[40]));
   AO22X1 U6526 (.IN1(\key_mem[11][41] ), .IN2(n6496), .IN3(\key_mem[6][41] ), .IN4(n6481)
          , .Q(n5847));
   AO221X1 U6527 (.IN1(\key_mem[4][41] ), .IN2(n6526), .IN3(\key_mem[5][41] ), .IN4(n6511)
          , .IN5(n5847), .Q(n5853));
   AO222X1 U6528 (.IN1(\key_mem[9][41] ), .IN2(n6571), .IN3(\key_mem[8][41] ), .IN4(n6556)
          , .IN5(\key_mem[10][41] ), .IN6(n6541), .Q(n5852));
   AO22X1 U6529 (.IN1(\key_mem[3][41] ), .IN2(n6601), .IN3(\key_mem[14][41] ), .IN4(n6586)
          , .Q(n5848));
   AO221X1 U6530 (.IN1(\key_mem[12][41] ), .IN2(n6631), .IN3(\key_mem[13][41] ), .IN4(
          n6616), .IN5(n5848), .Q(n5851));
   AO22X1 U6531 (.IN1(\key_mem[7][41] ), .IN2(n6661), .IN3(\key_mem[2][41] ), .IN4(n6646)
          , .Q(n5849));
   AO221X1 U6532 (.IN1(\key_mem[0][41] ), .IN2(n6691), .IN3(\key_mem[1][41] ), .IN4(n6676)
          , .IN5(n5849), .Q(n5850));
   OR4X1 U6533 (.IN1(n5853), .IN2(n5852), .IN3(n5851), .IN4(n5850), .Q(round_key[41]));
   AO22X1 U6534 (.IN1(\key_mem[11][42] ), .IN2(n6496), .IN3(\key_mem[6][42] ), .IN4(n6481)
          , .Q(n5854));
   AO221X1 U6535 (.IN1(\key_mem[4][42] ), .IN2(n6526), .IN3(\key_mem[5][42] ), .IN4(n6511)
          , .IN5(n5854), .Q(n5860));
   AO222X1 U6536 (.IN1(\key_mem[9][42] ), .IN2(n6571), .IN3(\key_mem[8][42] ), .IN4(n6556)
          , .IN5(\key_mem[10][42] ), .IN6(n6541), .Q(n5859));
   AO22X1 U6537 (.IN1(\key_mem[3][42] ), .IN2(n6601), .IN3(\key_mem[14][42] ), .IN4(n6586)
          , .Q(n5855));
   AO221X1 U6538 (.IN1(\key_mem[12][42] ), .IN2(n6631), .IN3(\key_mem[13][42] ), .IN4(
          n6616), .IN5(n5855), .Q(n5858));
   AO22X1 U6539 (.IN1(\key_mem[7][42] ), .IN2(n6661), .IN3(\key_mem[2][42] ), .IN4(n6646)
          , .Q(n5856));
   AO221X1 U6540 (.IN1(\key_mem[0][42] ), .IN2(n6691), .IN3(\key_mem[1][42] ), .IN4(n6676)
          , .IN5(n5856), .Q(n5857));
   OR4X1 U6541 (.IN1(n5860), .IN2(n5859), .IN3(n5858), .IN4(n5857), .Q(round_key[42]));
   AO22X1 U6542 (.IN1(\key_mem[11][43] ), .IN2(n6496), .IN3(\key_mem[6][43] ), .IN4(n6481)
          , .Q(n5861));
   AO221X1 U6543 (.IN1(\key_mem[4][43] ), .IN2(n6526), .IN3(\key_mem[5][43] ), .IN4(n6511)
          , .IN5(n5861), .Q(n5867));
   AO222X1 U6544 (.IN1(\key_mem[9][43] ), .IN2(n6571), .IN3(\key_mem[8][43] ), .IN4(n6556)
          , .IN5(\key_mem[10][43] ), .IN6(n6541), .Q(n5866));
   AO22X1 U6545 (.IN1(\key_mem[3][43] ), .IN2(n6601), .IN3(\key_mem[14][43] ), .IN4(n6586)
          , .Q(n5862));
   AO221X1 U6546 (.IN1(\key_mem[12][43] ), .IN2(n6631), .IN3(\key_mem[13][43] ), .IN4(
          n6616), .IN5(n5862), .Q(n5865));
   AO22X1 U6547 (.IN1(\key_mem[7][43] ), .IN2(n6661), .IN3(\key_mem[2][43] ), .IN4(n6646)
          , .Q(n5863));
   AO221X1 U6548 (.IN1(\key_mem[0][43] ), .IN2(n6691), .IN3(\key_mem[1][43] ), .IN4(n6676)
          , .IN5(n5863), .Q(n5864));
   OR4X1 U6549 (.IN1(n5867), .IN2(n5866), .IN3(n5865), .IN4(n5864), .Q(round_key[43]));
   AO22X1 U6550 (.IN1(\key_mem[11][44] ), .IN2(n6496), .IN3(\key_mem[6][44] ), .IN4(n6481)
          , .Q(n5868));
   AO221X1 U6551 (.IN1(\key_mem[4][44] ), .IN2(n6526), .IN3(\key_mem[5][44] ), .IN4(n6511)
          , .IN5(n5868), .Q(n5874));
   AO222X1 U6552 (.IN1(\key_mem[9][44] ), .IN2(n6571), .IN3(\key_mem[8][44] ), .IN4(n6556)
          , .IN5(\key_mem[10][44] ), .IN6(n6541), .Q(n5873));
   AO22X1 U6553 (.IN1(\key_mem[3][44] ), .IN2(n6601), .IN3(\key_mem[14][44] ), .IN4(n6586)
          , .Q(n5869));
   AO221X1 U6554 (.IN1(\key_mem[12][44] ), .IN2(n6631), .IN3(\key_mem[13][44] ), .IN4(
          n6616), .IN5(n5869), .Q(n5872));
   AO22X1 U6555 (.IN1(\key_mem[7][44] ), .IN2(n6661), .IN3(\key_mem[2][44] ), .IN4(n6646)
          , .Q(n5870));
   AO221X1 U6556 (.IN1(\key_mem[0][44] ), .IN2(n6691), .IN3(\key_mem[1][44] ), .IN4(n6676)
          , .IN5(n5870), .Q(n5871));
   OR4X1 U6557 (.IN1(n5874), .IN2(n5873), .IN3(n5872), .IN4(n5871), .Q(round_key[44]));
   AO22X1 U6558 (.IN1(\key_mem[11][45] ), .IN2(n6496), .IN3(\key_mem[6][45] ), .IN4(n6481)
          , .Q(n5875));
   AO221X1 U6559 (.IN1(\key_mem[4][45] ), .IN2(n6526), .IN3(\key_mem[5][45] ), .IN4(n6511)
          , .IN5(n5875), .Q(n5881));
   AO222X1 U6560 (.IN1(\key_mem[9][45] ), .IN2(n6571), .IN3(\key_mem[8][45] ), .IN4(n6556)
          , .IN5(\key_mem[10][45] ), .IN6(n6541), .Q(n5880));
   AO22X1 U6561 (.IN1(\key_mem[3][45] ), .IN2(n6601), .IN3(\key_mem[14][45] ), .IN4(n6586)
          , .Q(n5876));
   AO221X1 U6562 (.IN1(\key_mem[12][45] ), .IN2(n6631), .IN3(\key_mem[13][45] ), .IN4(
          n6616), .IN5(n5876), .Q(n5879));
   AO22X1 U6563 (.IN1(\key_mem[7][45] ), .IN2(n6661), .IN3(\key_mem[2][45] ), .IN4(n6646)
          , .Q(n5877));
   AO221X1 U6564 (.IN1(\key_mem[0][45] ), .IN2(n6691), .IN3(\key_mem[1][45] ), .IN4(n6676)
          , .IN5(n5877), .Q(n5878));
   OR4X1 U6565 (.IN1(n5881), .IN2(n5880), .IN3(n5879), .IN4(n5878), .Q(round_key[45]));
   AO22X1 U6566 (.IN1(\key_mem[11][46] ), .IN2(n6496), .IN3(\key_mem[6][46] ), .IN4(n6481)
          , .Q(n5882));
   AO221X1 U6567 (.IN1(\key_mem[4][46] ), .IN2(n6526), .IN3(\key_mem[5][46] ), .IN4(n6511)
          , .IN5(n5882), .Q(n5888));
   AO222X1 U6568 (.IN1(\key_mem[9][46] ), .IN2(n6571), .IN3(\key_mem[8][46] ), .IN4(n6556)
          , .IN5(\key_mem[10][46] ), .IN6(n6541), .Q(n5887));
   AO22X1 U6569 (.IN1(\key_mem[3][46] ), .IN2(n6601), .IN3(\key_mem[14][46] ), .IN4(n6586)
          , .Q(n5883));
   AO221X1 U6570 (.IN1(\key_mem[12][46] ), .IN2(n6631), .IN3(\key_mem[13][46] ), .IN4(
          n6616), .IN5(n5883), .Q(n5886));
   AO22X1 U6571 (.IN1(\key_mem[7][46] ), .IN2(n6661), .IN3(\key_mem[2][46] ), .IN4(n6646)
          , .Q(n5884));
   AO221X1 U6572 (.IN1(\key_mem[0][46] ), .IN2(n6691), .IN3(\key_mem[1][46] ), .IN4(n6676)
          , .IN5(n5884), .Q(n5885));
   OR4X1 U6573 (.IN1(n5888), .IN2(n5887), .IN3(n5886), .IN4(n5885), .Q(round_key[46]));
   AO22X1 U6574 (.IN1(\key_mem[11][47] ), .IN2(n6496), .IN3(\key_mem[6][47] ), .IN4(n6481)
          , .Q(n5889));
   AO221X1 U6575 (.IN1(\key_mem[4][47] ), .IN2(n6526), .IN3(\key_mem[5][47] ), .IN4(n6511)
          , .IN5(n5889), .Q(n5895));
   AO222X1 U6576 (.IN1(\key_mem[9][47] ), .IN2(n6571), .IN3(\key_mem[8][47] ), .IN4(n6556)
          , .IN5(\key_mem[10][47] ), .IN6(n6541), .Q(n5894));
   AO22X1 U6577 (.IN1(\key_mem[3][47] ), .IN2(n6601), .IN3(\key_mem[14][47] ), .IN4(n6586)
          , .Q(n5890));
   AO221X1 U6578 (.IN1(\key_mem[12][47] ), .IN2(n6631), .IN3(\key_mem[13][47] ), .IN4(
          n6616), .IN5(n5890), .Q(n5893));
   AO22X1 U6579 (.IN1(\key_mem[7][47] ), .IN2(n6661), .IN3(\key_mem[2][47] ), .IN4(n6646)
          , .Q(n5891));
   AO221X1 U6580 (.IN1(\key_mem[0][47] ), .IN2(n6691), .IN3(\key_mem[1][47] ), .IN4(n6676)
          , .IN5(n5891), .Q(n5892));
   OR4X1 U6581 (.IN1(n5895), .IN2(n5894), .IN3(n5893), .IN4(n5892), .Q(round_key[47]));
   AO22X1 U6582 (.IN1(\key_mem[11][48] ), .IN2(n6495), .IN3(\key_mem[6][48] ), .IN4(n6480)
          , .Q(n5896));
   AO221X1 U6583 (.IN1(\key_mem[4][48] ), .IN2(n6525), .IN3(\key_mem[5][48] ), .IN4(n6510)
          , .IN5(n5896), .Q(n5902));
   AO222X1 U6584 (.IN1(\key_mem[9][48] ), .IN2(n6570), .IN3(\key_mem[8][48] ), .IN4(n6555)
          , .IN5(\key_mem[10][48] ), .IN6(n6540), .Q(n5901));
   AO22X1 U6585 (.IN1(\key_mem[3][48] ), .IN2(n6600), .IN3(\key_mem[14][48] ), .IN4(n6585)
          , .Q(n5897));
   AO221X1 U6586 (.IN1(\key_mem[12][48] ), .IN2(n6630), .IN3(\key_mem[13][48] ), .IN4(
          n6615), .IN5(n5897), .Q(n5900));
   AO22X1 U6587 (.IN1(\key_mem[7][48] ), .IN2(n6660), .IN3(\key_mem[2][48] ), .IN4(n6645)
          , .Q(n5898));
   AO221X1 U6588 (.IN1(\key_mem[0][48] ), .IN2(n6690), .IN3(\key_mem[1][48] ), .IN4(n6675)
          , .IN5(n5898), .Q(n5899));
   OR4X1 U6589 (.IN1(n5902), .IN2(n5901), .IN3(n5900), .IN4(n5899), .Q(round_key[48]));
   AO22X1 U6590 (.IN1(\key_mem[11][49] ), .IN2(n6495), .IN3(\key_mem[6][49] ), .IN4(n6480)
          , .Q(n5903));
   AO221X1 U6591 (.IN1(\key_mem[4][49] ), .IN2(n6525), .IN3(\key_mem[5][49] ), .IN4(n6510)
          , .IN5(n5903), .Q(n5909));
   AO222X1 U6592 (.IN1(\key_mem[9][49] ), .IN2(n6570), .IN3(\key_mem[8][49] ), .IN4(n6555)
          , .IN5(\key_mem[10][49] ), .IN6(n6540), .Q(n5908));
   AO22X1 U6593 (.IN1(\key_mem[3][49] ), .IN2(n6600), .IN3(\key_mem[14][49] ), .IN4(n6585)
          , .Q(n5904));
   AO221X1 U6594 (.IN1(\key_mem[12][49] ), .IN2(n6630), .IN3(\key_mem[13][49] ), .IN4(
          n6615), .IN5(n5904), .Q(n5907));
   AO22X1 U6595 (.IN1(\key_mem[7][49] ), .IN2(n6660), .IN3(\key_mem[2][49] ), .IN4(n6645)
          , .Q(n5905));
   AO221X1 U6596 (.IN1(\key_mem[0][49] ), .IN2(n6690), .IN3(\key_mem[1][49] ), .IN4(n6675)
          , .IN5(n5905), .Q(n5906));
   OR4X1 U6597 (.IN1(n5909), .IN2(n5908), .IN3(n5907), .IN4(n5906), .Q(round_key[49]));
   AO22X1 U6598 (.IN1(\key_mem[11][50] ), .IN2(n6495), .IN3(\key_mem[6][50] ), .IN4(n6480)
          , .Q(n5910));
   AO221X1 U6599 (.IN1(\key_mem[4][50] ), .IN2(n6525), .IN3(\key_mem[5][50] ), .IN4(n6510)
          , .IN5(n5910), .Q(n5916));
   AO222X1 U6600 (.IN1(\key_mem[9][50] ), .IN2(n6570), .IN3(\key_mem[8][50] ), .IN4(n6555)
          , .IN5(\key_mem[10][50] ), .IN6(n6540), .Q(n5915));
   AO22X1 U6601 (.IN1(\key_mem[3][50] ), .IN2(n6600), .IN3(\key_mem[14][50] ), .IN4(n6585)
          , .Q(n5911));
   AO221X1 U6602 (.IN1(\key_mem[12][50] ), .IN2(n6630), .IN3(\key_mem[13][50] ), .IN4(
          n6615), .IN5(n5911), .Q(n5914));
   AO22X1 U6603 (.IN1(\key_mem[7][50] ), .IN2(n6660), .IN3(\key_mem[2][50] ), .IN4(n6645)
          , .Q(n5912));
   AO221X1 U6604 (.IN1(\key_mem[0][50] ), .IN2(n6690), .IN3(\key_mem[1][50] ), .IN4(n6675)
          , .IN5(n5912), .Q(n5913));
   OR4X1 U6605 (.IN1(n5916), .IN2(n5915), .IN3(n5914), .IN4(n5913), .Q(round_key[50]));
   AO22X1 U6606 (.IN1(\key_mem[11][51] ), .IN2(n6495), .IN3(\key_mem[6][51] ), .IN4(n6480)
          , .Q(n5917));
   AO221X1 U6607 (.IN1(\key_mem[4][51] ), .IN2(n6525), .IN3(\key_mem[5][51] ), .IN4(n6510)
          , .IN5(n5917), .Q(n5923));
   AO222X1 U6608 (.IN1(\key_mem[9][51] ), .IN2(n6570), .IN3(\key_mem[8][51] ), .IN4(n6555)
          , .IN5(\key_mem[10][51] ), .IN6(n6540), .Q(n5922));
   AO22X1 U6609 (.IN1(\key_mem[3][51] ), .IN2(n6600), .IN3(\key_mem[14][51] ), .IN4(n6585)
          , .Q(n5918));
   AO221X1 U6610 (.IN1(\key_mem[12][51] ), .IN2(n6630), .IN3(\key_mem[13][51] ), .IN4(
          n6615), .IN5(n5918), .Q(n5921));
   AO22X1 U6611 (.IN1(\key_mem[7][51] ), .IN2(n6660), .IN3(\key_mem[2][51] ), .IN4(n6645)
          , .Q(n5919));
   AO221X1 U6612 (.IN1(\key_mem[0][51] ), .IN2(n6690), .IN3(\key_mem[1][51] ), .IN4(n6675)
          , .IN5(n5919), .Q(n5920));
   OR4X1 U6613 (.IN1(n5923), .IN2(n5922), .IN3(n5921), .IN4(n5920), .Q(round_key[51]));
   AO22X1 U6614 (.IN1(\key_mem[11][52] ), .IN2(n6495), .IN3(\key_mem[6][52] ), .IN4(n6480)
          , .Q(n5924));
   AO221X1 U6615 (.IN1(\key_mem[4][52] ), .IN2(n6525), .IN3(\key_mem[5][52] ), .IN4(n6510)
          , .IN5(n5924), .Q(n5930));
   AO222X1 U6616 (.IN1(\key_mem[9][52] ), .IN2(n6570), .IN3(\key_mem[8][52] ), .IN4(n6555)
          , .IN5(\key_mem[10][52] ), .IN6(n6540), .Q(n5929));
   AO22X1 U6617 (.IN1(\key_mem[3][52] ), .IN2(n6600), .IN3(\key_mem[14][52] ), .IN4(n6585)
          , .Q(n5925));
   AO221X1 U6618 (.IN1(\key_mem[12][52] ), .IN2(n6630), .IN3(\key_mem[13][52] ), .IN4(
          n6615), .IN5(n5925), .Q(n5928));
   AO22X1 U6619 (.IN1(\key_mem[7][52] ), .IN2(n6660), .IN3(\key_mem[2][52] ), .IN4(n6645)
          , .Q(n5926));
   AO221X1 U6620 (.IN1(\key_mem[0][52] ), .IN2(n6690), .IN3(\key_mem[1][52] ), .IN4(n6675)
          , .IN5(n5926), .Q(n5927));
   OR4X1 U6621 (.IN1(n5930), .IN2(n5929), .IN3(n5928), .IN4(n5927), .Q(round_key[52]));
   AO22X1 U6622 (.IN1(\key_mem[11][53] ), .IN2(n6495), .IN3(\key_mem[6][53] ), .IN4(n6480)
          , .Q(n5931));
   AO221X1 U6623 (.IN1(\key_mem[4][53] ), .IN2(n6525), .IN3(\key_mem[5][53] ), .IN4(n6510)
          , .IN5(n5931), .Q(n5937));
   AO222X1 U6624 (.IN1(\key_mem[9][53] ), .IN2(n6570), .IN3(\key_mem[8][53] ), .IN4(n6555)
          , .IN5(\key_mem[10][53] ), .IN6(n6540), .Q(n5936));
   AO22X1 U6625 (.IN1(\key_mem[3][53] ), .IN2(n6600), .IN3(\key_mem[14][53] ), .IN4(n6585)
          , .Q(n5932));
   AO221X1 U6626 (.IN1(\key_mem[12][53] ), .IN2(n6630), .IN3(\key_mem[13][53] ), .IN4(
          n6615), .IN5(n5932), .Q(n5935));
   AO22X1 U6627 (.IN1(\key_mem[7][53] ), .IN2(n6660), .IN3(\key_mem[2][53] ), .IN4(n6645)
          , .Q(n5933));
   AO221X1 U6628 (.IN1(\key_mem[0][53] ), .IN2(n6690), .IN3(\key_mem[1][53] ), .IN4(n6675)
          , .IN5(n5933), .Q(n5934));
   OR4X1 U6629 (.IN1(n5937), .IN2(n5936), .IN3(n5935), .IN4(n5934), .Q(round_key[53]));
   AO22X1 U6630 (.IN1(\key_mem[11][54] ), .IN2(n6495), .IN3(\key_mem[6][54] ), .IN4(n6480)
          , .Q(n5938));
   AO221X1 U6631 (.IN1(\key_mem[4][54] ), .IN2(n6525), .IN3(\key_mem[5][54] ), .IN4(n6510)
          , .IN5(n5938), .Q(n5944));
   AO222X1 U6632 (.IN1(\key_mem[9][54] ), .IN2(n6570), .IN3(\key_mem[8][54] ), .IN4(n6555)
          , .IN5(\key_mem[10][54] ), .IN6(n6540), .Q(n5943));
   AO22X1 U6633 (.IN1(\key_mem[3][54] ), .IN2(n6600), .IN3(\key_mem[14][54] ), .IN4(n6585)
          , .Q(n5939));
   AO221X1 U6634 (.IN1(\key_mem[12][54] ), .IN2(n6630), .IN3(\key_mem[13][54] ), .IN4(
          n6615), .IN5(n5939), .Q(n5942));
   AO22X1 U6635 (.IN1(\key_mem[7][54] ), .IN2(n6660), .IN3(\key_mem[2][54] ), .IN4(n6645)
          , .Q(n5940));
   AO221X1 U6636 (.IN1(\key_mem[0][54] ), .IN2(n6690), .IN3(\key_mem[1][54] ), .IN4(n6675)
          , .IN5(n5940), .Q(n5941));
   OR4X1 U6637 (.IN1(n5944), .IN2(n5943), .IN3(n5942), .IN4(n5941), .Q(round_key[54]));
   AO22X1 U6638 (.IN1(\key_mem[11][55] ), .IN2(n6495), .IN3(\key_mem[6][55] ), .IN4(n6480)
          , .Q(n5945));
   AO221X1 U6639 (.IN1(\key_mem[4][55] ), .IN2(n6525), .IN3(\key_mem[5][55] ), .IN4(n6510)
          , .IN5(n5945), .Q(n5951));
   AO222X1 U6640 (.IN1(\key_mem[9][55] ), .IN2(n6570), .IN3(\key_mem[8][55] ), .IN4(n6555)
          , .IN5(\key_mem[10][55] ), .IN6(n6540), .Q(n5950));
   AO22X1 U6641 (.IN1(\key_mem[3][55] ), .IN2(n6600), .IN3(\key_mem[14][55] ), .IN4(n6585)
          , .Q(n5946));
   AO221X1 U6642 (.IN1(\key_mem[12][55] ), .IN2(n6630), .IN3(\key_mem[13][55] ), .IN4(
          n6615), .IN5(n5946), .Q(n5949));
   AO22X1 U6643 (.IN1(\key_mem[7][55] ), .IN2(n6660), .IN3(\key_mem[2][55] ), .IN4(n6645)
          , .Q(n5947));
   AO221X1 U6644 (.IN1(\key_mem[0][55] ), .IN2(n6690), .IN3(\key_mem[1][55] ), .IN4(n6675)
          , .IN5(n5947), .Q(n5948));
   OR4X1 U6645 (.IN1(n5951), .IN2(n5950), .IN3(n5949), .IN4(n5948), .Q(round_key[55]));
   AO22X1 U6646 (.IN1(\key_mem[11][56] ), .IN2(n6495), .IN3(\key_mem[6][56] ), .IN4(n6480)
          , .Q(n5952));
   AO221X1 U6647 (.IN1(\key_mem[4][56] ), .IN2(n6525), .IN3(\key_mem[5][56] ), .IN4(n6510)
          , .IN5(n5952), .Q(n5958));
   AO222X1 U6648 (.IN1(\key_mem[9][56] ), .IN2(n6570), .IN3(\key_mem[8][56] ), .IN4(n6555)
          , .IN5(\key_mem[10][56] ), .IN6(n6540), .Q(n5957));
   AO22X1 U6649 (.IN1(\key_mem[3][56] ), .IN2(n6600), .IN3(\key_mem[14][56] ), .IN4(n6585)
          , .Q(n5953));
   AO221X1 U6650 (.IN1(\key_mem[12][56] ), .IN2(n6630), .IN3(\key_mem[13][56] ), .IN4(
          n6615), .IN5(n5953), .Q(n5956));
   AO22X1 U6651 (.IN1(\key_mem[7][56] ), .IN2(n6660), .IN3(\key_mem[2][56] ), .IN4(n6645)
          , .Q(n5954));
   AO221X1 U6652 (.IN1(\key_mem[0][56] ), .IN2(n6690), .IN3(\key_mem[1][56] ), .IN4(n6675)
          , .IN5(n5954), .Q(n5955));
   OR4X1 U6653 (.IN1(n5958), .IN2(n5957), .IN3(n5956), .IN4(n5955), .Q(round_key[56]));
   AO22X1 U6654 (.IN1(\key_mem[11][57] ), .IN2(n6495), .IN3(\key_mem[6][57] ), .IN4(n6480)
          , .Q(n5959));
   AO221X1 U6655 (.IN1(\key_mem[4][57] ), .IN2(n6525), .IN3(\key_mem[5][57] ), .IN4(n6510)
          , .IN5(n5959), .Q(n5965));
   AO222X1 U6656 (.IN1(\key_mem[9][57] ), .IN2(n6570), .IN3(\key_mem[8][57] ), .IN4(n6555)
          , .IN5(\key_mem[10][57] ), .IN6(n6540), .Q(n5964));
   AO22X1 U6657 (.IN1(\key_mem[3][57] ), .IN2(n6600), .IN3(\key_mem[14][57] ), .IN4(n6585)
          , .Q(n5960));
   AO221X1 U6658 (.IN1(\key_mem[12][57] ), .IN2(n6630), .IN3(\key_mem[13][57] ), .IN4(
          n6615), .IN5(n5960), .Q(n5963));
   AO22X1 U6659 (.IN1(\key_mem[7][57] ), .IN2(n6660), .IN3(\key_mem[2][57] ), .IN4(n6645)
          , .Q(n5961));
   AO221X1 U6660 (.IN1(\key_mem[0][57] ), .IN2(n6690), .IN3(\key_mem[1][57] ), .IN4(n6675)
          , .IN5(n5961), .Q(n5962));
   OR4X1 U6661 (.IN1(n5965), .IN2(n5964), .IN3(n5963), .IN4(n5962), .Q(round_key[57]));
   AO22X1 U6662 (.IN1(\key_mem[11][58] ), .IN2(n6495), .IN3(\key_mem[6][58] ), .IN4(n6480)
          , .Q(n5966));
   AO221X1 U6663 (.IN1(\key_mem[4][58] ), .IN2(n6525), .IN3(\key_mem[5][58] ), .IN4(n6510)
          , .IN5(n5966), .Q(n5972));
   AO222X1 U6664 (.IN1(\key_mem[9][58] ), .IN2(n6570), .IN3(\key_mem[8][58] ), .IN4(n6555)
          , .IN5(\key_mem[10][58] ), .IN6(n6540), .Q(n5971));
   AO22X1 U6665 (.IN1(\key_mem[3][58] ), .IN2(n6600), .IN3(\key_mem[14][58] ), .IN4(n6585)
          , .Q(n5967));
   AO221X1 U6666 (.IN1(\key_mem[12][58] ), .IN2(n6630), .IN3(\key_mem[13][58] ), .IN4(
          n6615), .IN5(n5967), .Q(n5970));
   AO22X1 U6667 (.IN1(\key_mem[7][58] ), .IN2(n6660), .IN3(\key_mem[2][58] ), .IN4(n6645)
          , .Q(n5968));
   AO221X1 U6668 (.IN1(\key_mem[0][58] ), .IN2(n6690), .IN3(\key_mem[1][58] ), .IN4(n6675)
          , .IN5(n5968), .Q(n5969));
   OR4X1 U6669 (.IN1(n5972), .IN2(n5971), .IN3(n5970), .IN4(n5969), .Q(round_key[58]));
   AO22X1 U6670 (.IN1(\key_mem[11][59] ), .IN2(n6495), .IN3(\key_mem[6][59] ), .IN4(n6480)
          , .Q(n5973));
   AO221X1 U6671 (.IN1(\key_mem[4][59] ), .IN2(n6525), .IN3(\key_mem[5][59] ), .IN4(n6510)
          , .IN5(n5973), .Q(n5979));
   AO222X1 U6672 (.IN1(\key_mem[9][59] ), .IN2(n6570), .IN3(\key_mem[8][59] ), .IN4(n6555)
          , .IN5(\key_mem[10][59] ), .IN6(n6540), .Q(n5978));
   AO22X1 U6673 (.IN1(\key_mem[3][59] ), .IN2(n6600), .IN3(\key_mem[14][59] ), .IN4(n6585)
          , .Q(n5974));
   AO221X1 U6674 (.IN1(\key_mem[12][59] ), .IN2(n6630), .IN3(\key_mem[13][59] ), .IN4(
          n6615), .IN5(n5974), .Q(n5977));
   AO22X1 U6675 (.IN1(\key_mem[7][59] ), .IN2(n6660), .IN3(\key_mem[2][59] ), .IN4(n6645)
          , .Q(n5975));
   AO221X1 U6676 (.IN1(\key_mem[0][59] ), .IN2(n6690), .IN3(\key_mem[1][59] ), .IN4(n6675)
          , .IN5(n5975), .Q(n5976));
   OR4X1 U6677 (.IN1(n5979), .IN2(n5978), .IN3(n5977), .IN4(n5976), .Q(round_key[59]));
   AO22X1 U6678 (.IN1(\key_mem[11][60] ), .IN2(n6494), .IN3(\key_mem[6][60] ), .IN4(n6479)
          , .Q(n5980));
   AO221X1 U6679 (.IN1(\key_mem[4][60] ), .IN2(n6524), .IN3(\key_mem[5][60] ), .IN4(n6509)
          , .IN5(n5980), .Q(n5986));
   AO222X1 U6680 (.IN1(\key_mem[9][60] ), .IN2(n6569), .IN3(\key_mem[8][60] ), .IN4(n6554)
          , .IN5(\key_mem[10][60] ), .IN6(n6539), .Q(n5985));
   AO22X1 U6681 (.IN1(\key_mem[3][60] ), .IN2(n6599), .IN3(\key_mem[14][60] ), .IN4(n6584)
          , .Q(n5981));
   AO221X1 U6682 (.IN1(\key_mem[12][60] ), .IN2(n6629), .IN3(\key_mem[13][60] ), .IN4(
          n6614), .IN5(n5981), .Q(n5984));
   AO22X1 U6683 (.IN1(\key_mem[7][60] ), .IN2(n6659), .IN3(\key_mem[2][60] ), .IN4(n6644)
          , .Q(n5982));
   AO221X1 U6684 (.IN1(\key_mem[0][60] ), .IN2(n6689), .IN3(\key_mem[1][60] ), .IN4(n6674)
          , .IN5(n5982), .Q(n5983));
   OR4X1 U6685 (.IN1(n5986), .IN2(n5985), .IN3(n5984), .IN4(n5983), .Q(round_key[60]));
   AO22X1 U6686 (.IN1(\key_mem[11][61] ), .IN2(n6494), .IN3(\key_mem[6][61] ), .IN4(n6479)
          , .Q(n5987));
   AO221X1 U6687 (.IN1(\key_mem[4][61] ), .IN2(n6524), .IN3(\key_mem[5][61] ), .IN4(n6509)
          , .IN5(n5987), .Q(n5993));
   AO222X1 U6688 (.IN1(\key_mem[9][61] ), .IN2(n6569), .IN3(\key_mem[8][61] ), .IN4(n6554)
          , .IN5(\key_mem[10][61] ), .IN6(n6539), .Q(n5992));
   AO22X1 U6689 (.IN1(\key_mem[3][61] ), .IN2(n6599), .IN3(\key_mem[14][61] ), .IN4(n6584)
          , .Q(n5988));
   AO221X1 U6690 (.IN1(\key_mem[12][61] ), .IN2(n6629), .IN3(\key_mem[13][61] ), .IN4(
          n6614), .IN5(n5988), .Q(n5991));
   AO22X1 U6691 (.IN1(\key_mem[7][61] ), .IN2(n6659), .IN3(\key_mem[2][61] ), .IN4(n6644)
          , .Q(n5989));
   AO221X1 U6692 (.IN1(\key_mem[0][61] ), .IN2(n6689), .IN3(\key_mem[1][61] ), .IN4(n6674)
          , .IN5(n5989), .Q(n5990));
   OR4X1 U6693 (.IN1(n5993), .IN2(n5992), .IN3(n5991), .IN4(n5990), .Q(round_key[61]));
   AO22X1 U6694 (.IN1(\key_mem[11][62] ), .IN2(n6494), .IN3(\key_mem[6][62] ), .IN4(n6479)
          , .Q(n5994));
   AO221X1 U6695 (.IN1(\key_mem[4][62] ), .IN2(n6524), .IN3(\key_mem[5][62] ), .IN4(n6509)
          , .IN5(n5994), .Q(n6000));
   AO222X1 U6696 (.IN1(\key_mem[9][62] ), .IN2(n6569), .IN3(\key_mem[8][62] ), .IN4(n6554)
          , .IN5(\key_mem[10][62] ), .IN6(n6539), .Q(n5999));
   AO22X1 U6697 (.IN1(\key_mem[3][62] ), .IN2(n6599), .IN3(\key_mem[14][62] ), .IN4(n6584)
          , .Q(n5995));
   AO221X1 U6698 (.IN1(\key_mem[12][62] ), .IN2(n6629), .IN3(\key_mem[13][62] ), .IN4(
          n6614), .IN5(n5995), .Q(n5998));
   AO22X1 U6699 (.IN1(\key_mem[7][62] ), .IN2(n6659), .IN3(\key_mem[2][62] ), .IN4(n6644)
          , .Q(n5996));
   AO221X1 U6700 (.IN1(\key_mem[0][62] ), .IN2(n6689), .IN3(\key_mem[1][62] ), .IN4(n6674)
          , .IN5(n5996), .Q(n5997));
   OR4X1 U6701 (.IN1(n6000), .IN2(n5999), .IN3(n5998), .IN4(n5997), .Q(round_key[62]));
   AO22X1 U6702 (.IN1(\key_mem[11][63] ), .IN2(n6494), .IN3(\key_mem[6][63] ), .IN4(n6479)
          , .Q(n6001));
   AO221X1 U6703 (.IN1(\key_mem[4][63] ), .IN2(n6524), .IN3(\key_mem[5][63] ), .IN4(n6509)
          , .IN5(n6001), .Q(n6007));
   AO222X1 U6704 (.IN1(\key_mem[9][63] ), .IN2(n6569), .IN3(\key_mem[8][63] ), .IN4(n6554)
          , .IN5(\key_mem[10][63] ), .IN6(n6539), .Q(n6006));
   AO22X1 U6705 (.IN1(\key_mem[3][63] ), .IN2(n6599), .IN3(\key_mem[14][63] ), .IN4(n6584)
          , .Q(n6002));
   AO221X1 U6706 (.IN1(\key_mem[12][63] ), .IN2(n6629), .IN3(\key_mem[13][63] ), .IN4(
          n6614), .IN5(n6002), .Q(n6005));
   AO22X1 U6707 (.IN1(\key_mem[7][63] ), .IN2(n6659), .IN3(\key_mem[2][63] ), .IN4(n6644)
          , .Q(n6003));
   AO221X1 U6708 (.IN1(\key_mem[0][63] ), .IN2(n6689), .IN3(\key_mem[1][63] ), .IN4(n6674)
          , .IN5(n6003), .Q(n6004));
   OR4X1 U6709 (.IN1(n6007), .IN2(n6006), .IN3(n6005), .IN4(n6004), .Q(round_key[63]));
   AO22X1 U6710 (.IN1(\key_mem[11][64] ), .IN2(n6494), .IN3(\key_mem[6][64] ), .IN4(n6479)
          , .Q(n6008));
   AO221X1 U6711 (.IN1(\key_mem[4][64] ), .IN2(n6524), .IN3(\key_mem[5][64] ), .IN4(n6509)
          , .IN5(n6008), .Q(n6014));
   AO222X1 U6712 (.IN1(\key_mem[9][64] ), .IN2(n6569), .IN3(\key_mem[8][64] ), .IN4(n6554)
          , .IN5(\key_mem[10][64] ), .IN6(n6539), .Q(n6013));
   AO22X1 U6713 (.IN1(\key_mem[3][64] ), .IN2(n6599), .IN3(\key_mem[14][64] ), .IN4(n6584)
          , .Q(n6009));
   AO221X1 U6714 (.IN1(\key_mem[12][64] ), .IN2(n6629), .IN3(\key_mem[13][64] ), .IN4(
          n6614), .IN5(n6009), .Q(n6012));
   AO22X1 U6715 (.IN1(\key_mem[7][64] ), .IN2(n6659), .IN3(\key_mem[2][64] ), .IN4(n6644)
          , .Q(n6010));
   AO221X1 U6716 (.IN1(\key_mem[0][64] ), .IN2(n6689), .IN3(\key_mem[1][64] ), .IN4(n6674)
          , .IN5(n6010), .Q(n6011));
   OR4X1 U6717 (.IN1(n6014), .IN2(n6013), .IN3(n6012), .IN4(n6011), .Q(round_key[64]));
   AO22X1 U6718 (.IN1(\key_mem[11][65] ), .IN2(n6494), .IN3(\key_mem[6][65] ), .IN4(n6479)
          , .Q(n6015));
   AO221X1 U6719 (.IN1(\key_mem[4][65] ), .IN2(n6524), .IN3(\key_mem[5][65] ), .IN4(n6509)
          , .IN5(n6015), .Q(n6021));
   AO222X1 U6720 (.IN1(\key_mem[9][65] ), .IN2(n6569), .IN3(\key_mem[8][65] ), .IN4(n6554)
          , .IN5(\key_mem[10][65] ), .IN6(n6539), .Q(n6020));
   AO22X1 U6721 (.IN1(\key_mem[3][65] ), .IN2(n6599), .IN3(\key_mem[14][65] ), .IN4(n6584)
          , .Q(n6016));
   AO221X1 U6722 (.IN1(\key_mem[12][65] ), .IN2(n6629), .IN3(\key_mem[13][65] ), .IN4(
          n6614), .IN5(n6016), .Q(n6019));
   AO22X1 U6723 (.IN1(\key_mem[7][65] ), .IN2(n6659), .IN3(\key_mem[2][65] ), .IN4(n6644)
          , .Q(n6017));
   AO221X1 U6724 (.IN1(\key_mem[0][65] ), .IN2(n6689), .IN3(\key_mem[1][65] ), .IN4(n6674)
          , .IN5(n6017), .Q(n6018));
   OR4X1 U6725 (.IN1(n6021), .IN2(n6020), .IN3(n6019), .IN4(n6018), .Q(round_key[65]));
   AO22X1 U6726 (.IN1(\key_mem[11][66] ), .IN2(n6494), .IN3(\key_mem[6][66] ), .IN4(n6479)
          , .Q(n6022));
   AO221X1 U6727 (.IN1(\key_mem[4][66] ), .IN2(n6524), .IN3(\key_mem[5][66] ), .IN4(n6509)
          , .IN5(n6022), .Q(n6028));
   AO222X1 U6728 (.IN1(\key_mem[9][66] ), .IN2(n6569), .IN3(\key_mem[8][66] ), .IN4(n6554)
          , .IN5(\key_mem[10][66] ), .IN6(n6539), .Q(n6027));
   AO22X1 U6729 (.IN1(\key_mem[3][66] ), .IN2(n6599), .IN3(\key_mem[14][66] ), .IN4(n6584)
          , .Q(n6023));
   AO221X1 U6730 (.IN1(\key_mem[12][66] ), .IN2(n6629), .IN3(\key_mem[13][66] ), .IN4(
          n6614), .IN5(n6023), .Q(n6026));
   AO22X1 U6731 (.IN1(\key_mem[7][66] ), .IN2(n6659), .IN3(\key_mem[2][66] ), .IN4(n6644)
          , .Q(n6024));
   AO221X1 U6732 (.IN1(\key_mem[0][66] ), .IN2(n6689), .IN3(\key_mem[1][66] ), .IN4(n6674)
          , .IN5(n6024), .Q(n6025));
   OR4X1 U6733 (.IN1(n6028), .IN2(n6027), .IN3(n6026), .IN4(n6025), .Q(round_key[66]));
   AO22X1 U6734 (.IN1(\key_mem[11][67] ), .IN2(n6494), .IN3(\key_mem[6][67] ), .IN4(n6479)
          , .Q(n6029));
   AO221X1 U6735 (.IN1(\key_mem[4][67] ), .IN2(n6524), .IN3(\key_mem[5][67] ), .IN4(n6509)
          , .IN5(n6029), .Q(n6035));
   AO222X1 U6736 (.IN1(\key_mem[9][67] ), .IN2(n6569), .IN3(\key_mem[8][67] ), .IN4(n6554)
          , .IN5(\key_mem[10][67] ), .IN6(n6539), .Q(n6034));
   AO22X1 U6737 (.IN1(\key_mem[3][67] ), .IN2(n6599), .IN3(\key_mem[14][67] ), .IN4(n6584)
          , .Q(n6030));
   AO221X1 U6738 (.IN1(\key_mem[12][67] ), .IN2(n6629), .IN3(\key_mem[13][67] ), .IN4(
          n6614), .IN5(n6030), .Q(n6033));
   AO22X1 U6739 (.IN1(\key_mem[7][67] ), .IN2(n6659), .IN3(\key_mem[2][67] ), .IN4(n6644)
          , .Q(n6031));
   AO221X1 U6740 (.IN1(\key_mem[0][67] ), .IN2(n6689), .IN3(\key_mem[1][67] ), .IN4(n6674)
          , .IN5(n6031), .Q(n6032));
   OR4X1 U6741 (.IN1(n6035), .IN2(n6034), .IN3(n6033), .IN4(n6032), .Q(round_key[67]));
   AO22X1 U6742 (.IN1(\key_mem[11][68] ), .IN2(n6494), .IN3(\key_mem[6][68] ), .IN4(n6479)
          , .Q(n6036));
   AO221X1 U6743 (.IN1(\key_mem[4][68] ), .IN2(n6524), .IN3(\key_mem[5][68] ), .IN4(n6509)
          , .IN5(n6036), .Q(n6042));
   AO222X1 U6744 (.IN1(\key_mem[9][68] ), .IN2(n6569), .IN3(\key_mem[8][68] ), .IN4(n6554)
          , .IN5(\key_mem[10][68] ), .IN6(n6539), .Q(n6041));
   AO22X1 U6745 (.IN1(\key_mem[3][68] ), .IN2(n6599), .IN3(\key_mem[14][68] ), .IN4(n6584)
          , .Q(n6037));
   AO221X1 U6746 (.IN1(\key_mem[12][68] ), .IN2(n6629), .IN3(\key_mem[13][68] ), .IN4(
          n6614), .IN5(n6037), .Q(n6040));
   AO22X1 U6747 (.IN1(\key_mem[7][68] ), .IN2(n6659), .IN3(\key_mem[2][68] ), .IN4(n6644)
          , .Q(n6038));
   AO221X1 U6748 (.IN1(\key_mem[0][68] ), .IN2(n6689), .IN3(\key_mem[1][68] ), .IN4(n6674)
          , .IN5(n6038), .Q(n6039));
   OR4X1 U6749 (.IN1(n6042), .IN2(n6041), .IN3(n6040), .IN4(n6039), .Q(round_key[68]));
   AO22X1 U6750 (.IN1(\key_mem[11][69] ), .IN2(n6494), .IN3(\key_mem[6][69] ), .IN4(n6479)
          , .Q(n6043));
   AO221X1 U6751 (.IN1(\key_mem[4][69] ), .IN2(n6524), .IN3(\key_mem[5][69] ), .IN4(n6509)
          , .IN5(n6043), .Q(n6049));
   AO222X1 U6752 (.IN1(\key_mem[9][69] ), .IN2(n6569), .IN3(\key_mem[8][69] ), .IN4(n6554)
          , .IN5(\key_mem[10][69] ), .IN6(n6539), .Q(n6048));
   AO22X1 U6753 (.IN1(\key_mem[3][69] ), .IN2(n6599), .IN3(\key_mem[14][69] ), .IN4(n6584)
          , .Q(n6044));
   AO221X1 U6754 (.IN1(\key_mem[12][69] ), .IN2(n6629), .IN3(\key_mem[13][69] ), .IN4(
          n6614), .IN5(n6044), .Q(n6047));
   AO22X1 U6755 (.IN1(\key_mem[7][69] ), .IN2(n6659), .IN3(\key_mem[2][69] ), .IN4(n6644)
          , .Q(n6045));
   AO221X1 U6756 (.IN1(\key_mem[0][69] ), .IN2(n6689), .IN3(\key_mem[1][69] ), .IN4(n6674)
          , .IN5(n6045), .Q(n6046));
   OR4X1 U6757 (.IN1(n6049), .IN2(n6048), .IN3(n6047), .IN4(n6046), .Q(round_key[69]));
   AO22X1 U6758 (.IN1(\key_mem[11][70] ), .IN2(n6494), .IN3(\key_mem[6][70] ), .IN4(n6479)
          , .Q(n6050));
   AO221X1 U6759 (.IN1(\key_mem[4][70] ), .IN2(n6524), .IN3(\key_mem[5][70] ), .IN4(n6509)
          , .IN5(n6050), .Q(n6056));
   AO222X1 U6760 (.IN1(\key_mem[9][70] ), .IN2(n6569), .IN3(\key_mem[8][70] ), .IN4(n6554)
          , .IN5(\key_mem[10][70] ), .IN6(n6539), .Q(n6055));
   AO22X1 U6761 (.IN1(\key_mem[3][70] ), .IN2(n6599), .IN3(\key_mem[14][70] ), .IN4(n6584)
          , .Q(n6051));
   AO221X1 U6762 (.IN1(\key_mem[12][70] ), .IN2(n6629), .IN3(\key_mem[13][70] ), .IN4(
          n6614), .IN5(n6051), .Q(n6054));
   AO22X1 U6763 (.IN1(\key_mem[7][70] ), .IN2(n6659), .IN3(\key_mem[2][70] ), .IN4(n6644)
          , .Q(n6052));
   AO221X1 U6764 (.IN1(\key_mem[0][70] ), .IN2(n6689), .IN3(\key_mem[1][70] ), .IN4(n6674)
          , .IN5(n6052), .Q(n6053));
   OR4X1 U6765 (.IN1(n6056), .IN2(n6055), .IN3(n6054), .IN4(n6053), .Q(round_key[70]));
   AO22X1 U6766 (.IN1(\key_mem[11][71] ), .IN2(n6494), .IN3(\key_mem[6][71] ), .IN4(n6479)
          , .Q(n6057));
   AO221X1 U6767 (.IN1(\key_mem[4][71] ), .IN2(n6524), .IN3(\key_mem[5][71] ), .IN4(n6509)
          , .IN5(n6057), .Q(n6063));
   AO222X1 U6768 (.IN1(\key_mem[9][71] ), .IN2(n6569), .IN3(\key_mem[8][71] ), .IN4(n6554)
          , .IN5(\key_mem[10][71] ), .IN6(n6539), .Q(n6062));
   AO22X1 U6769 (.IN1(\key_mem[3][71] ), .IN2(n6599), .IN3(\key_mem[14][71] ), .IN4(n6584)
          , .Q(n6058));
   AO221X1 U6770 (.IN1(\key_mem[12][71] ), .IN2(n6629), .IN3(\key_mem[13][71] ), .IN4(
          n6614), .IN5(n6058), .Q(n6061));
   AO22X1 U6771 (.IN1(\key_mem[7][71] ), .IN2(n6659), .IN3(\key_mem[2][71] ), .IN4(n6644)
          , .Q(n6059));
   AO221X1 U6772 (.IN1(\key_mem[0][71] ), .IN2(n6689), .IN3(\key_mem[1][71] ), .IN4(n6674)
          , .IN5(n6059), .Q(n6060));
   OR4X1 U6773 (.IN1(n6063), .IN2(n6062), .IN3(n6061), .IN4(n6060), .Q(round_key[71]));
   AO22X1 U6774 (.IN1(\key_mem[11][72] ), .IN2(n6493), .IN3(\key_mem[6][72] ), .IN4(n6478)
          , .Q(n6064));
   AO221X1 U6775 (.IN1(\key_mem[4][72] ), .IN2(n6523), .IN3(\key_mem[5][72] ), .IN4(n6508)
          , .IN5(n6064), .Q(n6070));
   AO222X1 U6776 (.IN1(\key_mem[9][72] ), .IN2(n6568), .IN3(\key_mem[8][72] ), .IN4(n6553)
          , .IN5(\key_mem[10][72] ), .IN6(n6538), .Q(n6069));
   AO22X1 U6777 (.IN1(\key_mem[3][72] ), .IN2(n6598), .IN3(\key_mem[14][72] ), .IN4(n6583)
          , .Q(n6065));
   AO221X1 U6778 (.IN1(\key_mem[12][72] ), .IN2(n6628), .IN3(\key_mem[13][72] ), .IN4(
          n6613), .IN5(n6065), .Q(n6068));
   AO22X1 U6779 (.IN1(\key_mem[7][72] ), .IN2(n6658), .IN3(\key_mem[2][72] ), .IN4(n6643)
          , .Q(n6066));
   AO221X1 U6780 (.IN1(\key_mem[0][72] ), .IN2(n6688), .IN3(\key_mem[1][72] ), .IN4(n6673)
          , .IN5(n6066), .Q(n6067));
   OR4X1 U6781 (.IN1(n6070), .IN2(n6069), .IN3(n6068), .IN4(n6067), .Q(round_key[72]));
   AO22X1 U6782 (.IN1(\key_mem[11][73] ), .IN2(n6493), .IN3(\key_mem[6][73] ), .IN4(n6478)
          , .Q(n6071));
   AO221X1 U6783 (.IN1(\key_mem[4][73] ), .IN2(n6523), .IN3(\key_mem[5][73] ), .IN4(n6508)
          , .IN5(n6071), .Q(n6077));
   AO222X1 U6784 (.IN1(\key_mem[9][73] ), .IN2(n6568), .IN3(\key_mem[8][73] ), .IN4(n6553)
          , .IN5(\key_mem[10][73] ), .IN6(n6538), .Q(n6076));
   AO22X1 U6785 (.IN1(\key_mem[3][73] ), .IN2(n6598), .IN3(\key_mem[14][73] ), .IN4(n6583)
          , .Q(n6072));
   AO221X1 U6786 (.IN1(\key_mem[12][73] ), .IN2(n6628), .IN3(\key_mem[13][73] ), .IN4(
          n6613), .IN5(n6072), .Q(n6075));
   AO22X1 U6787 (.IN1(\key_mem[7][73] ), .IN2(n6658), .IN3(\key_mem[2][73] ), .IN4(n6643)
          , .Q(n6073));
   AO221X1 U6788 (.IN1(\key_mem[0][73] ), .IN2(n6688), .IN3(\key_mem[1][73] ), .IN4(n6673)
          , .IN5(n6073), .Q(n6074));
   OR4X1 U6789 (.IN1(n6077), .IN2(n6076), .IN3(n6075), .IN4(n6074), .Q(round_key[73]));
   AO22X1 U6790 (.IN1(\key_mem[11][74] ), .IN2(n6493), .IN3(\key_mem[6][74] ), .IN4(n6478)
          , .Q(n6078));
   AO221X1 U6791 (.IN1(\key_mem[4][74] ), .IN2(n6523), .IN3(\key_mem[5][74] ), .IN4(n6508)
          , .IN5(n6078), .Q(n6084));
   AO222X1 U6792 (.IN1(\key_mem[9][74] ), .IN2(n6568), .IN3(\key_mem[8][74] ), .IN4(n6553)
          , .IN5(\key_mem[10][74] ), .IN6(n6538), .Q(n6083));
   AO22X1 U6793 (.IN1(\key_mem[3][74] ), .IN2(n6598), .IN3(\key_mem[14][74] ), .IN4(n6583)
          , .Q(n6079));
   AO221X1 U6794 (.IN1(\key_mem[12][74] ), .IN2(n6628), .IN3(\key_mem[13][74] ), .IN4(
          n6613), .IN5(n6079), .Q(n6082));
   AO22X1 U6795 (.IN1(\key_mem[7][74] ), .IN2(n6658), .IN3(\key_mem[2][74] ), .IN4(n6643)
          , .Q(n6080));
   AO221X1 U6796 (.IN1(\key_mem[0][74] ), .IN2(n6688), .IN3(\key_mem[1][74] ), .IN4(n6673)
          , .IN5(n6080), .Q(n6081));
   OR4X1 U6797 (.IN1(n6084), .IN2(n6083), .IN3(n6082), .IN4(n6081), .Q(round_key[74]));
   AO22X1 U6798 (.IN1(\key_mem[11][75] ), .IN2(n6493), .IN3(\key_mem[6][75] ), .IN4(n6478)
          , .Q(n6085));
   AO221X1 U6799 (.IN1(\key_mem[4][75] ), .IN2(n6523), .IN3(\key_mem[5][75] ), .IN4(n6508)
          , .IN5(n6085), .Q(n6091));
   AO222X1 U6800 (.IN1(\key_mem[9][75] ), .IN2(n6568), .IN3(\key_mem[8][75] ), .IN4(n6553)
          , .IN5(\key_mem[10][75] ), .IN6(n6538), .Q(n6090));
   AO22X1 U6801 (.IN1(\key_mem[3][75] ), .IN2(n6598), .IN3(\key_mem[14][75] ), .IN4(n6583)
          , .Q(n6086));
   AO221X1 U6802 (.IN1(\key_mem[12][75] ), .IN2(n6628), .IN3(\key_mem[13][75] ), .IN4(
          n6613), .IN5(n6086), .Q(n6089));
   AO22X1 U6803 (.IN1(\key_mem[7][75] ), .IN2(n6658), .IN3(\key_mem[2][75] ), .IN4(n6643)
          , .Q(n6087));
   AO221X1 U6804 (.IN1(\key_mem[0][75] ), .IN2(n6688), .IN3(\key_mem[1][75] ), .IN4(n6673)
          , .IN5(n6087), .Q(n6088));
   OR4X1 U6805 (.IN1(n6091), .IN2(n6090), .IN3(n6089), .IN4(n6088), .Q(round_key[75]));
   AO22X1 U6806 (.IN1(\key_mem[11][76] ), .IN2(n6493), .IN3(\key_mem[6][76] ), .IN4(n6478)
          , .Q(n6092));
   AO221X1 U6807 (.IN1(\key_mem[4][76] ), .IN2(n6523), .IN3(\key_mem[5][76] ), .IN4(n6508)
          , .IN5(n6092), .Q(n6098));
   AO222X1 U6808 (.IN1(\key_mem[9][76] ), .IN2(n6568), .IN3(\key_mem[8][76] ), .IN4(n6553)
          , .IN5(\key_mem[10][76] ), .IN6(n6538), .Q(n6097));
   AO22X1 U6809 (.IN1(\key_mem[3][76] ), .IN2(n6598), .IN3(\key_mem[14][76] ), .IN4(n6583)
          , .Q(n6093));
   AO221X1 U6810 (.IN1(\key_mem[12][76] ), .IN2(n6628), .IN3(\key_mem[13][76] ), .IN4(
          n6613), .IN5(n6093), .Q(n6096));
   AO22X1 U6811 (.IN1(\key_mem[7][76] ), .IN2(n6658), .IN3(\key_mem[2][76] ), .IN4(n6643)
          , .Q(n6094));
   AO221X1 U6812 (.IN1(\key_mem[0][76] ), .IN2(n6688), .IN3(\key_mem[1][76] ), .IN4(n6673)
          , .IN5(n6094), .Q(n6095));
   OR4X1 U6813 (.IN1(n6098), .IN2(n6097), .IN3(n6096), .IN4(n6095), .Q(round_key[76]));
   AO22X1 U6814 (.IN1(\key_mem[11][77] ), .IN2(n6493), .IN3(\key_mem[6][77] ), .IN4(n6478)
          , .Q(n6099));
   AO221X1 U6815 (.IN1(\key_mem[4][77] ), .IN2(n6523), .IN3(\key_mem[5][77] ), .IN4(n6508)
          , .IN5(n6099), .Q(n6105));
   AO222X1 U6816 (.IN1(\key_mem[9][77] ), .IN2(n6568), .IN3(\key_mem[8][77] ), .IN4(n6553)
          , .IN5(\key_mem[10][77] ), .IN6(n6538), .Q(n6104));
   AO22X1 U6817 (.IN1(\key_mem[3][77] ), .IN2(n6598), .IN3(\key_mem[14][77] ), .IN4(n6583)
          , .Q(n6100));
   AO221X1 U6818 (.IN1(\key_mem[12][77] ), .IN2(n6628), .IN3(\key_mem[13][77] ), .IN4(
          n6613), .IN5(n6100), .Q(n6103));
   AO22X1 U6819 (.IN1(\key_mem[7][77] ), .IN2(n6658), .IN3(\key_mem[2][77] ), .IN4(n6643)
          , .Q(n6101));
   AO221X1 U6820 (.IN1(\key_mem[0][77] ), .IN2(n6688), .IN3(\key_mem[1][77] ), .IN4(n6673)
          , .IN5(n6101), .Q(n6102));
   OR4X1 U6821 (.IN1(n6105), .IN2(n6104), .IN3(n6103), .IN4(n6102), .Q(round_key[77]));
   AO22X1 U6822 (.IN1(\key_mem[11][78] ), .IN2(n6493), .IN3(\key_mem[6][78] ), .IN4(n6478)
          , .Q(n6106));
   AO221X1 U6823 (.IN1(\key_mem[4][78] ), .IN2(n6523), .IN3(\key_mem[5][78] ), .IN4(n6508)
          , .IN5(n6106), .Q(n6112));
   AO222X1 U6824 (.IN1(\key_mem[9][78] ), .IN2(n6568), .IN3(\key_mem[8][78] ), .IN4(n6553)
          , .IN5(\key_mem[10][78] ), .IN6(n6538), .Q(n6111));
   AO22X1 U6825 (.IN1(\key_mem[3][78] ), .IN2(n6598), .IN3(\key_mem[14][78] ), .IN4(n6583)
          , .Q(n6107));
   AO221X1 U6826 (.IN1(\key_mem[12][78] ), .IN2(n6628), .IN3(\key_mem[13][78] ), .IN4(
          n6613), .IN5(n6107), .Q(n6110));
   AO22X1 U6827 (.IN1(\key_mem[7][78] ), .IN2(n6658), .IN3(\key_mem[2][78] ), .IN4(n6643)
          , .Q(n6108));
   AO221X1 U6828 (.IN1(\key_mem[0][78] ), .IN2(n6688), .IN3(\key_mem[1][78] ), .IN4(n6673)
          , .IN5(n6108), .Q(n6109));
   OR4X1 U6829 (.IN1(n6112), .IN2(n6111), .IN3(n6110), .IN4(n6109), .Q(round_key[78]));
   AO22X1 U6830 (.IN1(\key_mem[11][79] ), .IN2(n6493), .IN3(\key_mem[6][79] ), .IN4(n6478)
          , .Q(n6113));
   AO221X1 U6831 (.IN1(\key_mem[4][79] ), .IN2(n6523), .IN3(\key_mem[5][79] ), .IN4(n6508)
          , .IN5(n6113), .Q(n6119));
   AO222X1 U6832 (.IN1(\key_mem[9][79] ), .IN2(n6568), .IN3(\key_mem[8][79] ), .IN4(n6553)
          , .IN5(\key_mem[10][79] ), .IN6(n6538), .Q(n6118));
   AO22X1 U6833 (.IN1(\key_mem[3][79] ), .IN2(n6598), .IN3(\key_mem[14][79] ), .IN4(n6583)
          , .Q(n6114));
   AO221X1 U6834 (.IN1(\key_mem[12][79] ), .IN2(n6628), .IN3(\key_mem[13][79] ), .IN4(
          n6613), .IN5(n6114), .Q(n6117));
   AO22X1 U6835 (.IN1(\key_mem[7][79] ), .IN2(n6658), .IN3(\key_mem[2][79] ), .IN4(n6643)
          , .Q(n6115));
   AO221X1 U6836 (.IN1(\key_mem[0][79] ), .IN2(n6688), .IN3(\key_mem[1][79] ), .IN4(n6673)
          , .IN5(n6115), .Q(n6116));
   OR4X1 U6837 (.IN1(n6119), .IN2(n6118), .IN3(n6117), .IN4(n6116), .Q(round_key[79]));
   AO22X1 U6838 (.IN1(\key_mem[11][80] ), .IN2(n6493), .IN3(\key_mem[6][80] ), .IN4(n6478)
          , .Q(n6120));
   AO221X1 U6839 (.IN1(\key_mem[4][80] ), .IN2(n6523), .IN3(\key_mem[5][80] ), .IN4(n6508)
          , .IN5(n6120), .Q(n6126));
   AO222X1 U6840 (.IN1(\key_mem[9][80] ), .IN2(n6568), .IN3(\key_mem[8][80] ), .IN4(n6553)
          , .IN5(\key_mem[10][80] ), .IN6(n6538), .Q(n6125));
   AO22X1 U6841 (.IN1(\key_mem[3][80] ), .IN2(n6598), .IN3(\key_mem[14][80] ), .IN4(n6583)
          , .Q(n6121));
   AO221X1 U6842 (.IN1(\key_mem[12][80] ), .IN2(n6628), .IN3(\key_mem[13][80] ), .IN4(
          n6613), .IN5(n6121), .Q(n6124));
   AO22X1 U6843 (.IN1(\key_mem[7][80] ), .IN2(n6658), .IN3(\key_mem[2][80] ), .IN4(n6643)
          , .Q(n6122));
   AO221X1 U6844 (.IN1(\key_mem[0][80] ), .IN2(n6688), .IN3(\key_mem[1][80] ), .IN4(n6673)
          , .IN5(n6122), .Q(n6123));
   OR4X1 U6845 (.IN1(n6126), .IN2(n6125), .IN3(n6124), .IN4(n6123), .Q(round_key[80]));
   AO22X1 U6846 (.IN1(\key_mem[11][81] ), .IN2(n6493), .IN3(\key_mem[6][81] ), .IN4(n6478)
          , .Q(n6127));
   AO221X1 U6847 (.IN1(\key_mem[4][81] ), .IN2(n6523), .IN3(\key_mem[5][81] ), .IN4(n6508)
          , .IN5(n6127), .Q(n6133));
   AO222X1 U6848 (.IN1(\key_mem[9][81] ), .IN2(n6568), .IN3(\key_mem[8][81] ), .IN4(n6553)
          , .IN5(\key_mem[10][81] ), .IN6(n6538), .Q(n6132));
   AO22X1 U6849 (.IN1(\key_mem[3][81] ), .IN2(n6598), .IN3(\key_mem[14][81] ), .IN4(n6583)
          , .Q(n6128));
   AO221X1 U6850 (.IN1(\key_mem[12][81] ), .IN2(n6628), .IN3(\key_mem[13][81] ), .IN4(
          n6613), .IN5(n6128), .Q(n6131));
   AO22X1 U6851 (.IN1(\key_mem[7][81] ), .IN2(n6658), .IN3(\key_mem[2][81] ), .IN4(n6643)
          , .Q(n6129));
   AO221X1 U6852 (.IN1(\key_mem[0][81] ), .IN2(n6688), .IN3(\key_mem[1][81] ), .IN4(n6673)
          , .IN5(n6129), .Q(n6130));
   OR4X1 U6853 (.IN1(n6133), .IN2(n6132), .IN3(n6131), .IN4(n6130), .Q(round_key[81]));
   AO22X1 U6854 (.IN1(\key_mem[11][82] ), .IN2(n6493), .IN3(\key_mem[6][82] ), .IN4(n6478)
          , .Q(n6134));
   AO221X1 U6855 (.IN1(\key_mem[4][82] ), .IN2(n6523), .IN3(\key_mem[5][82] ), .IN4(n6508)
          , .IN5(n6134), .Q(n6140));
   AO222X1 U6856 (.IN1(\key_mem[9][82] ), .IN2(n6568), .IN3(\key_mem[8][82] ), .IN4(n6553)
          , .IN5(\key_mem[10][82] ), .IN6(n6538), .Q(n6139));
   AO22X1 U6857 (.IN1(\key_mem[3][82] ), .IN2(n6598), .IN3(\key_mem[14][82] ), .IN4(n6583)
          , .Q(n6135));
   AO221X1 U6858 (.IN1(\key_mem[12][82] ), .IN2(n6628), .IN3(\key_mem[13][82] ), .IN4(
          n6613), .IN5(n6135), .Q(n6138));
   AO22X1 U6859 (.IN1(\key_mem[7][82] ), .IN2(n6658), .IN3(\key_mem[2][82] ), .IN4(n6643)
          , .Q(n6136));
   AO221X1 U6860 (.IN1(\key_mem[0][82] ), .IN2(n6688), .IN3(\key_mem[1][82] ), .IN4(n6673)
          , .IN5(n6136), .Q(n6137));
   OR4X1 U6861 (.IN1(n6140), .IN2(n6139), .IN3(n6138), .IN4(n6137), .Q(round_key[82]));
   AO22X1 U6862 (.IN1(\key_mem[11][83] ), .IN2(n6493), .IN3(\key_mem[6][83] ), .IN4(n6478)
          , .Q(n6141));
   AO221X1 U6863 (.IN1(\key_mem[4][83] ), .IN2(n6523), .IN3(\key_mem[5][83] ), .IN4(n6508)
          , .IN5(n6141), .Q(n6147));
   AO222X1 U6864 (.IN1(\key_mem[9][83] ), .IN2(n6568), .IN3(\key_mem[8][83] ), .IN4(n6553)
          , .IN5(\key_mem[10][83] ), .IN6(n6538), .Q(n6146));
   AO22X1 U6865 (.IN1(\key_mem[3][83] ), .IN2(n6598), .IN3(\key_mem[14][83] ), .IN4(n6583)
          , .Q(n6142));
   AO221X1 U6866 (.IN1(\key_mem[12][83] ), .IN2(n6628), .IN3(\key_mem[13][83] ), .IN4(
          n6613), .IN5(n6142), .Q(n6145));
   AO22X1 U6867 (.IN1(\key_mem[7][83] ), .IN2(n6658), .IN3(\key_mem[2][83] ), .IN4(n6643)
          , .Q(n6143));
   AO221X1 U6868 (.IN1(\key_mem[0][83] ), .IN2(n6688), .IN3(\key_mem[1][83] ), .IN4(n6673)
          , .IN5(n6143), .Q(n6144));
   OR4X1 U6869 (.IN1(n6147), .IN2(n6146), .IN3(n6145), .IN4(n6144), .Q(round_key[83]));
   AO22X1 U6870 (.IN1(\key_mem[11][84] ), .IN2(n6492), .IN3(\key_mem[6][84] ), .IN4(n6477)
          , .Q(n6148));
   AO221X1 U6871 (.IN1(\key_mem[4][84] ), .IN2(n6522), .IN3(\key_mem[5][84] ), .IN4(n6507)
          , .IN5(n6148), .Q(n6154));
   AO222X1 U6872 (.IN1(\key_mem[9][84] ), .IN2(n6567), .IN3(\key_mem[8][84] ), .IN4(n6552)
          , .IN5(\key_mem[10][84] ), .IN6(n6537), .Q(n6153));
   AO22X1 U6873 (.IN1(\key_mem[3][84] ), .IN2(n6597), .IN3(\key_mem[14][84] ), .IN4(n6582)
          , .Q(n6149));
   AO221X1 U6874 (.IN1(\key_mem[12][84] ), .IN2(n6627), .IN3(\key_mem[13][84] ), .IN4(
          n6612), .IN5(n6149), .Q(n6152));
   AO22X1 U6875 (.IN1(\key_mem[7][84] ), .IN2(n6657), .IN3(\key_mem[2][84] ), .IN4(n6642)
          , .Q(n6150));
   AO221X1 U6876 (.IN1(\key_mem[0][84] ), .IN2(n6687), .IN3(\key_mem[1][84] ), .IN4(n6672)
          , .IN5(n6150), .Q(n6151));
   OR4X1 U6877 (.IN1(n6154), .IN2(n6153), .IN3(n6152), .IN4(n6151), .Q(round_key[84]));
   AO22X1 U6878 (.IN1(\key_mem[11][85] ), .IN2(n6492), .IN3(\key_mem[6][85] ), .IN4(n6477)
          , .Q(n6155));
   AO221X1 U6879 (.IN1(\key_mem[4][85] ), .IN2(n6522), .IN3(\key_mem[5][85] ), .IN4(n6507)
          , .IN5(n6155), .Q(n6161));
   AO222X1 U6880 (.IN1(\key_mem[9][85] ), .IN2(n6567), .IN3(\key_mem[8][85] ), .IN4(n6552)
          , .IN5(\key_mem[10][85] ), .IN6(n6537), .Q(n6160));
   AO22X1 U6881 (.IN1(\key_mem[3][85] ), .IN2(n6597), .IN3(\key_mem[14][85] ), .IN4(n6582)
          , .Q(n6156));
   AO221X1 U6882 (.IN1(\key_mem[12][85] ), .IN2(n6627), .IN3(\key_mem[13][85] ), .IN4(
          n6612), .IN5(n6156), .Q(n6159));
   AO22X1 U6883 (.IN1(\key_mem[7][85] ), .IN2(n6657), .IN3(\key_mem[2][85] ), .IN4(n6642)
          , .Q(n6157));
   AO221X1 U6884 (.IN1(\key_mem[0][85] ), .IN2(n6687), .IN3(\key_mem[1][85] ), .IN4(n6672)
          , .IN5(n6157), .Q(n6158));
   OR4X1 U6885 (.IN1(n6161), .IN2(n6160), .IN3(n6159), .IN4(n6158), .Q(round_key[85]));
   AO22X1 U6886 (.IN1(\key_mem[11][86] ), .IN2(n6492), .IN3(\key_mem[6][86] ), .IN4(n6477)
          , .Q(n6162));
   AO221X1 U6887 (.IN1(\key_mem[4][86] ), .IN2(n6522), .IN3(\key_mem[5][86] ), .IN4(n6507)
          , .IN5(n6162), .Q(n6168));
   AO222X1 U6888 (.IN1(\key_mem[9][86] ), .IN2(n6567), .IN3(\key_mem[8][86] ), .IN4(n6552)
          , .IN5(\key_mem[10][86] ), .IN6(n6537), .Q(n6167));
   AO22X1 U6889 (.IN1(\key_mem[3][86] ), .IN2(n6597), .IN3(\key_mem[14][86] ), .IN4(n6582)
          , .Q(n6163));
   AO221X1 U6890 (.IN1(\key_mem[12][86] ), .IN2(n6627), .IN3(\key_mem[13][86] ), .IN4(
          n6612), .IN5(n6163), .Q(n6166));
   AO22X1 U6891 (.IN1(\key_mem[7][86] ), .IN2(n6657), .IN3(\key_mem[2][86] ), .IN4(n6642)
          , .Q(n6164));
   AO221X1 U6892 (.IN1(\key_mem[0][86] ), .IN2(n6687), .IN3(\key_mem[1][86] ), .IN4(n6672)
          , .IN5(n6164), .Q(n6165));
   OR4X1 U6893 (.IN1(n6168), .IN2(n6167), .IN3(n6166), .IN4(n6165), .Q(round_key[86]));
   AO22X1 U6894 (.IN1(\key_mem[11][87] ), .IN2(n6492), .IN3(\key_mem[6][87] ), .IN4(n6477)
          , .Q(n6169));
   AO221X1 U6895 (.IN1(\key_mem[4][87] ), .IN2(n6522), .IN3(\key_mem[5][87] ), .IN4(n6507)
          , .IN5(n6169), .Q(n6175));
   AO222X1 U6896 (.IN1(\key_mem[9][87] ), .IN2(n6567), .IN3(\key_mem[8][87] ), .IN4(n6552)
          , .IN5(\key_mem[10][87] ), .IN6(n6537), .Q(n6174));
   AO22X1 U6897 (.IN1(\key_mem[3][87] ), .IN2(n6597), .IN3(\key_mem[14][87] ), .IN4(n6582)
          , .Q(n6170));
   AO221X1 U6898 (.IN1(\key_mem[12][87] ), .IN2(n6627), .IN3(\key_mem[13][87] ), .IN4(
          n6612), .IN5(n6170), .Q(n6173));
   AO22X1 U6899 (.IN1(\key_mem[7][87] ), .IN2(n6657), .IN3(\key_mem[2][87] ), .IN4(n6642)
          , .Q(n6171));
   AO221X1 U6900 (.IN1(\key_mem[0][87] ), .IN2(n6687), .IN3(\key_mem[1][87] ), .IN4(n6672)
          , .IN5(n6171), .Q(n6172));
   OR4X1 U6901 (.IN1(n6175), .IN2(n6174), .IN3(n6173), .IN4(n6172), .Q(round_key[87]));
   AO22X1 U6902 (.IN1(\key_mem[11][88] ), .IN2(n6492), .IN3(\key_mem[6][88] ), .IN4(n6477)
          , .Q(n6176));
   AO221X1 U6903 (.IN1(\key_mem[4][88] ), .IN2(n6522), .IN3(\key_mem[5][88] ), .IN4(n6507)
          , .IN5(n6176), .Q(n6182));
   AO222X1 U6904 (.IN1(\key_mem[9][88] ), .IN2(n6567), .IN3(\key_mem[8][88] ), .IN4(n6552)
          , .IN5(\key_mem[10][88] ), .IN6(n6537), .Q(n6181));
   AO22X1 U6905 (.IN1(\key_mem[3][88] ), .IN2(n6597), .IN3(\key_mem[14][88] ), .IN4(n6582)
          , .Q(n6177));
   AO221X1 U6906 (.IN1(\key_mem[12][88] ), .IN2(n6627), .IN3(\key_mem[13][88] ), .IN4(
          n6612), .IN5(n6177), .Q(n6180));
   AO22X1 U6907 (.IN1(\key_mem[7][88] ), .IN2(n6657), .IN3(\key_mem[2][88] ), .IN4(n6642)
          , .Q(n6178));
   AO221X1 U6908 (.IN1(\key_mem[0][88] ), .IN2(n6687), .IN3(\key_mem[1][88] ), .IN4(n6672)
          , .IN5(n6178), .Q(n6179));
   OR4X1 U6909 (.IN1(n6182), .IN2(n6181), .IN3(n6180), .IN4(n6179), .Q(round_key[88]));
   AO22X1 U6910 (.IN1(\key_mem[11][89] ), .IN2(n6492), .IN3(\key_mem[6][89] ), .IN4(n6477)
          , .Q(n6183));
   AO221X1 U6911 (.IN1(\key_mem[4][89] ), .IN2(n6522), .IN3(\key_mem[5][89] ), .IN4(n6507)
          , .IN5(n6183), .Q(n6189));
   AO222X1 U6912 (.IN1(\key_mem[9][89] ), .IN2(n6567), .IN3(\key_mem[8][89] ), .IN4(n6552)
          , .IN5(\key_mem[10][89] ), .IN6(n6537), .Q(n6188));
   AO22X1 U6913 (.IN1(\key_mem[3][89] ), .IN2(n6597), .IN3(\key_mem[14][89] ), .IN4(n6582)
          , .Q(n6184));
   AO221X1 U6914 (.IN1(\key_mem[12][89] ), .IN2(n6627), .IN3(\key_mem[13][89] ), .IN4(
          n6612), .IN5(n6184), .Q(n6187));
   AO22X1 U6915 (.IN1(\key_mem[7][89] ), .IN2(n6657), .IN3(\key_mem[2][89] ), .IN4(n6642)
          , .Q(n6185));
   AO221X1 U6916 (.IN1(\key_mem[0][89] ), .IN2(n6687), .IN3(\key_mem[1][89] ), .IN4(n6672)
          , .IN5(n6185), .Q(n6186));
   OR4X1 U6917 (.IN1(n6189), .IN2(n6188), .IN3(n6187), .IN4(n6186), .Q(round_key[89]));
   AO22X1 U6918 (.IN1(\key_mem[11][90] ), .IN2(n6492), .IN3(\key_mem[6][90] ), .IN4(n6477)
          , .Q(n6190));
   AO221X1 U6919 (.IN1(\key_mem[4][90] ), .IN2(n6522), .IN3(\key_mem[5][90] ), .IN4(n6507)
          , .IN5(n6190), .Q(n6196));
   AO222X1 U6920 (.IN1(\key_mem[9][90] ), .IN2(n6567), .IN3(\key_mem[8][90] ), .IN4(n6552)
          , .IN5(\key_mem[10][90] ), .IN6(n6537), .Q(n6195));
   AO22X1 U6921 (.IN1(\key_mem[3][90] ), .IN2(n6597), .IN3(\key_mem[14][90] ), .IN4(n6582)
          , .Q(n6191));
   AO221X1 U6922 (.IN1(\key_mem[12][90] ), .IN2(n6627), .IN3(\key_mem[13][90] ), .IN4(
          n6612), .IN5(n6191), .Q(n6194));
   AO22X1 U6923 (.IN1(\key_mem[7][90] ), .IN2(n6657), .IN3(\key_mem[2][90] ), .IN4(n6642)
          , .Q(n6192));
   AO221X1 U6924 (.IN1(\key_mem[0][90] ), .IN2(n6687), .IN3(\key_mem[1][90] ), .IN4(n6672)
          , .IN5(n6192), .Q(n6193));
   OR4X1 U6925 (.IN1(n6196), .IN2(n6195), .IN3(n6194), .IN4(n6193), .Q(round_key[90]));
   AO22X1 U6926 (.IN1(\key_mem[11][91] ), .IN2(n6492), .IN3(\key_mem[6][91] ), .IN4(n6477)
          , .Q(n6197));
   AO221X1 U6927 (.IN1(\key_mem[4][91] ), .IN2(n6522), .IN3(\key_mem[5][91] ), .IN4(n6507)
          , .IN5(n6197), .Q(n6203));
   AO222X1 U6928 (.IN1(\key_mem[9][91] ), .IN2(n6567), .IN3(\key_mem[8][91] ), .IN4(n6552)
          , .IN5(\key_mem[10][91] ), .IN6(n6537), .Q(n6202));
   AO22X1 U6929 (.IN1(\key_mem[3][91] ), .IN2(n6597), .IN3(\key_mem[14][91] ), .IN4(n6582)
          , .Q(n6198));
   AO221X1 U6930 (.IN1(\key_mem[12][91] ), .IN2(n6627), .IN3(\key_mem[13][91] ), .IN4(
          n6612), .IN5(n6198), .Q(n6201));
   AO22X1 U6931 (.IN1(\key_mem[7][91] ), .IN2(n6657), .IN3(\key_mem[2][91] ), .IN4(n6642)
          , .Q(n6199));
   AO221X1 U6932 (.IN1(\key_mem[0][91] ), .IN2(n6687), .IN3(\key_mem[1][91] ), .IN4(n6672)
          , .IN5(n6199), .Q(n6200));
   OR4X1 U6933 (.IN1(n6203), .IN2(n6202), .IN3(n6201), .IN4(n6200), .Q(round_key[91]));
   AO22X1 U6934 (.IN1(\key_mem[11][92] ), .IN2(n6492), .IN3(\key_mem[6][92] ), .IN4(n6477)
          , .Q(n6204));
   AO221X1 U6935 (.IN1(\key_mem[4][92] ), .IN2(n6522), .IN3(\key_mem[5][92] ), .IN4(n6507)
          , .IN5(n6204), .Q(n6210));
   AO222X1 U6936 (.IN1(\key_mem[9][92] ), .IN2(n6567), .IN3(\key_mem[8][92] ), .IN4(n6552)
          , .IN5(\key_mem[10][92] ), .IN6(n6537), .Q(n6209));
   AO22X1 U6937 (.IN1(\key_mem[3][92] ), .IN2(n6597), .IN3(\key_mem[14][92] ), .IN4(n6582)
          , .Q(n6205));
   AO221X1 U6938 (.IN1(\key_mem[12][92] ), .IN2(n6627), .IN3(\key_mem[13][92] ), .IN4(
          n6612), .IN5(n6205), .Q(n6208));
   AO22X1 U6939 (.IN1(\key_mem[7][92] ), .IN2(n6657), .IN3(\key_mem[2][92] ), .IN4(n6642)
          , .Q(n6206));
   AO221X1 U6940 (.IN1(\key_mem[0][92] ), .IN2(n6687), .IN3(\key_mem[1][92] ), .IN4(n6672)
          , .IN5(n6206), .Q(n6207));
   OR4X1 U6941 (.IN1(n6210), .IN2(n6209), .IN3(n6208), .IN4(n6207), .Q(round_key[92]));
   AO22X1 U6942 (.IN1(\key_mem[11][93] ), .IN2(n6492), .IN3(\key_mem[6][93] ), .IN4(n6477)
          , .Q(n6211));
   AO221X1 U6943 (.IN1(\key_mem[4][93] ), .IN2(n6522), .IN3(\key_mem[5][93] ), .IN4(n6507)
          , .IN5(n6211), .Q(n6217));
   AO222X1 U6944 (.IN1(\key_mem[9][93] ), .IN2(n6567), .IN3(\key_mem[8][93] ), .IN4(n6552)
          , .IN5(\key_mem[10][93] ), .IN6(n6537), .Q(n6216));
   AO22X1 U6945 (.IN1(\key_mem[3][93] ), .IN2(n6597), .IN3(\key_mem[14][93] ), .IN4(n6582)
          , .Q(n6212));
   AO221X1 U6946 (.IN1(\key_mem[12][93] ), .IN2(n6627), .IN3(\key_mem[13][93] ), .IN4(
          n6612), .IN5(n6212), .Q(n6215));
   AO22X1 U6947 (.IN1(\key_mem[7][93] ), .IN2(n6657), .IN3(\key_mem[2][93] ), .IN4(n6642)
          , .Q(n6213));
   AO221X1 U6948 (.IN1(\key_mem[0][93] ), .IN2(n6687), .IN3(\key_mem[1][93] ), .IN4(n6672)
          , .IN5(n6213), .Q(n6214));
   OR4X1 U6949 (.IN1(n6217), .IN2(n6216), .IN3(n6215), .IN4(n6214), .Q(round_key[93]));
   AO22X1 U6950 (.IN1(\key_mem[11][94] ), .IN2(n6492), .IN3(\key_mem[6][94] ), .IN4(n6477)
          , .Q(n6218));
   AO221X1 U6951 (.IN1(\key_mem[4][94] ), .IN2(n6522), .IN3(\key_mem[5][94] ), .IN4(n6507)
          , .IN5(n6218), .Q(n6224));
   AO222X1 U6952 (.IN1(\key_mem[9][94] ), .IN2(n6567), .IN3(\key_mem[8][94] ), .IN4(n6552)
          , .IN5(\key_mem[10][94] ), .IN6(n6537), .Q(n6223));
   AO22X1 U6953 (.IN1(\key_mem[3][94] ), .IN2(n6597), .IN3(\key_mem[14][94] ), .IN4(n6582)
          , .Q(n6219));
   AO221X1 U6954 (.IN1(\key_mem[12][94] ), .IN2(n6627), .IN3(\key_mem[13][94] ), .IN4(
          n6612), .IN5(n6219), .Q(n6222));
   AO22X1 U6955 (.IN1(\key_mem[7][94] ), .IN2(n6657), .IN3(\key_mem[2][94] ), .IN4(n6642)
          , .Q(n6220));
   AO221X1 U6956 (.IN1(\key_mem[0][94] ), .IN2(n6687), .IN3(\key_mem[1][94] ), .IN4(n6672)
          , .IN5(n6220), .Q(n6221));
   OR4X1 U6957 (.IN1(n6224), .IN2(n6223), .IN3(n6222), .IN4(n6221), .Q(round_key[94]));
   AO22X1 U6958 (.IN1(\key_mem[11][95] ), .IN2(n6492), .IN3(\key_mem[6][95] ), .IN4(n6477)
          , .Q(n6225));
   AO221X1 U6959 (.IN1(\key_mem[4][95] ), .IN2(n6522), .IN3(\key_mem[5][95] ), .IN4(n6507)
          , .IN5(n6225), .Q(n6231));
   AO222X1 U6960 (.IN1(\key_mem[9][95] ), .IN2(n6567), .IN3(\key_mem[8][95] ), .IN4(n6552)
          , .IN5(\key_mem[10][95] ), .IN6(n6537), .Q(n6230));
   AO22X1 U6961 (.IN1(\key_mem[3][95] ), .IN2(n6597), .IN3(\key_mem[14][95] ), .IN4(n6582)
          , .Q(n6226));
   AO221X1 U6962 (.IN1(\key_mem[12][95] ), .IN2(n6627), .IN3(\key_mem[13][95] ), .IN4(
          n6612), .IN5(n6226), .Q(n6229));
   AO22X1 U6963 (.IN1(\key_mem[7][95] ), .IN2(n6657), .IN3(\key_mem[2][95] ), .IN4(n6642)
          , .Q(n6227));
   AO221X1 U6964 (.IN1(\key_mem[0][95] ), .IN2(n6687), .IN3(\key_mem[1][95] ), .IN4(n6672)
          , .IN5(n6227), .Q(n6228));
   OR4X1 U6965 (.IN1(n6231), .IN2(n6230), .IN3(n6229), .IN4(n6228), .Q(round_key[95]));
   AO22X1 U6966 (.IN1(\key_mem[11][96] ), .IN2(n6491), .IN3(\key_mem[6][96] ), .IN4(n6476)
          , .Q(n6232));
   AO221X1 U6967 (.IN1(\key_mem[4][96] ), .IN2(n6521), .IN3(\key_mem[5][96] ), .IN4(n6506)
          , .IN5(n6232), .Q(n6238));
   AO222X1 U6968 (.IN1(\key_mem[9][96] ), .IN2(n6566), .IN3(\key_mem[8][96] ), .IN4(n6551)
          , .IN5(\key_mem[10][96] ), .IN6(n6536), .Q(n6237));
   AO22X1 U6969 (.IN1(\key_mem[3][96] ), .IN2(n6596), .IN3(\key_mem[14][96] ), .IN4(n6581)
          , .Q(n6233));
   AO221X1 U6970 (.IN1(\key_mem[12][96] ), .IN2(n6626), .IN3(\key_mem[13][96] ), .IN4(
          n6611), .IN5(n6233), .Q(n6236));
   AO22X1 U6971 (.IN1(\key_mem[7][96] ), .IN2(n6656), .IN3(\key_mem[2][96] ), .IN4(n6641)
          , .Q(n6234));
   AO221X1 U6972 (.IN1(\key_mem[0][96] ), .IN2(n6686), .IN3(\key_mem[1][96] ), .IN4(n6671)
          , .IN5(n6234), .Q(n6235));
   OR4X1 U6973 (.IN1(n6238), .IN2(n6237), .IN3(n6236), .IN4(n6235), .Q(round_key[96]));
   AO22X1 U6974 (.IN1(\key_mem[11][97] ), .IN2(n6491), .IN3(\key_mem[6][97] ), .IN4(n6476)
          , .Q(n6239));
   AO221X1 U6975 (.IN1(\key_mem[4][97] ), .IN2(n6521), .IN3(\key_mem[5][97] ), .IN4(n6506)
          , .IN5(n6239), .Q(n6245));
   AO222X1 U6976 (.IN1(\key_mem[9][97] ), .IN2(n6566), .IN3(\key_mem[8][97] ), .IN4(n6551)
          , .IN5(\key_mem[10][97] ), .IN6(n6536), .Q(n6244));
   AO22X1 U6977 (.IN1(\key_mem[3][97] ), .IN2(n6596), .IN3(\key_mem[14][97] ), .IN4(n6581)
          , .Q(n6240));
   AO221X1 U6978 (.IN1(\key_mem[12][97] ), .IN2(n6626), .IN3(\key_mem[13][97] ), .IN4(
          n6611), .IN5(n6240), .Q(n6243));
   AO22X1 U6979 (.IN1(\key_mem[7][97] ), .IN2(n6656), .IN3(\key_mem[2][97] ), .IN4(n6641)
          , .Q(n6241));
   AO221X1 U6980 (.IN1(\key_mem[0][97] ), .IN2(n6686), .IN3(\key_mem[1][97] ), .IN4(n6671)
          , .IN5(n6241), .Q(n6242));
   OR4X1 U6981 (.IN1(n6245), .IN2(n6244), .IN3(n6243), .IN4(n6242), .Q(round_key[97]));
   AO22X1 U6982 (.IN1(\key_mem[11][98] ), .IN2(n6491), .IN3(\key_mem[6][98] ), .IN4(n6476)
          , .Q(n6246));
   AO221X1 U6983 (.IN1(\key_mem[4][98] ), .IN2(n6521), .IN3(\key_mem[5][98] ), .IN4(n6506)
          , .IN5(n6246), .Q(n6252));
   AO222X1 U6984 (.IN1(\key_mem[9][98] ), .IN2(n6566), .IN3(\key_mem[8][98] ), .IN4(n6551)
          , .IN5(\key_mem[10][98] ), .IN6(n6536), .Q(n6251));
   AO22X1 U6985 (.IN1(\key_mem[3][98] ), .IN2(n6596), .IN3(\key_mem[14][98] ), .IN4(n6581)
          , .Q(n6247));
   AO221X1 U6986 (.IN1(\key_mem[12][98] ), .IN2(n6626), .IN3(\key_mem[13][98] ), .IN4(
          n6611), .IN5(n6247), .Q(n6250));
   AO22X1 U6987 (.IN1(\key_mem[7][98] ), .IN2(n6656), .IN3(\key_mem[2][98] ), .IN4(n6641)
          , .Q(n6248));
   AO221X1 U6988 (.IN1(\key_mem[0][98] ), .IN2(n6686), .IN3(\key_mem[1][98] ), .IN4(n6671)
          , .IN5(n6248), .Q(n6249));
   OR4X1 U6989 (.IN1(n6252), .IN2(n6251), .IN3(n6250), .IN4(n6249), .Q(round_key[98]));
   AO22X1 U6990 (.IN1(\key_mem[11][99] ), .IN2(n6491), .IN3(\key_mem[6][99] ), .IN4(n6476)
          , .Q(n6253));
   AO221X1 U6991 (.IN1(\key_mem[4][99] ), .IN2(n6521), .IN3(\key_mem[5][99] ), .IN4(n6506)
          , .IN5(n6253), .Q(n6259));
   AO222X1 U6992 (.IN1(\key_mem[9][99] ), .IN2(n6566), .IN3(\key_mem[8][99] ), .IN4(n6551)
          , .IN5(\key_mem[10][99] ), .IN6(n6536), .Q(n6258));
   AO22X1 U6993 (.IN1(\key_mem[3][99] ), .IN2(n6596), .IN3(\key_mem[14][99] ), .IN4(n6581)
          , .Q(n6254));
   AO221X1 U6994 (.IN1(\key_mem[12][99] ), .IN2(n6626), .IN3(\key_mem[13][99] ), .IN4(
          n6611), .IN5(n6254), .Q(n6257));
   AO22X1 U6995 (.IN1(\key_mem[7][99] ), .IN2(n6656), .IN3(\key_mem[2][99] ), .IN4(n6641)
          , .Q(n6255));
   AO221X1 U6996 (.IN1(\key_mem[0][99] ), .IN2(n6686), .IN3(\key_mem[1][99] ), .IN4(n6671)
          , .IN5(n6255), .Q(n6256));
   OR4X1 U6997 (.IN1(n6259), .IN2(n6258), .IN3(n6257), .IN4(n6256), .Q(round_key[99]));
   AO22X1 U6998 (.IN1(\key_mem[11][100] ), .IN2(n6491), .IN3(\key_mem[6][100] ), .IN4(
          n6476), .Q(n6260));
   AO221X1 U6999 (.IN1(\key_mem[4][100] ), .IN2(n6521), .IN3(\key_mem[5][100] ), .IN4(
          n6506), .IN5(n6260), .Q(n6266));
   AO222X1 U7000 (.IN1(\key_mem[9][100] ), .IN2(n6566), .IN3(\key_mem[8][100] ), .IN4(
          n6551), .IN5(\key_mem[10][100] ), .IN6(n6536), .Q(n6265));
   AO22X1 U7001 (.IN1(\key_mem[3][100] ), .IN2(n6596), .IN3(\key_mem[14][100] ), .IN4(
          n6581), .Q(n6261));
   AO221X1 U7002 (.IN1(\key_mem[12][100] ), .IN2(n6626), .IN3(\key_mem[13][100] ), .IN4(
          n6611), .IN5(n6261), .Q(n6264));
   AO22X1 U7003 (.IN1(\key_mem[7][100] ), .IN2(n6656), .IN3(\key_mem[2][100] ), .IN4(n6641)
          , .Q(n6262));
   AO221X1 U7004 (.IN1(\key_mem[0][100] ), .IN2(n6686), .IN3(\key_mem[1][100] ), .IN4(
          n6671), .IN5(n6262), .Q(n6263));
   OR4X1 U7005 (.IN1(n6266), .IN2(n6265), .IN3(n6264), .IN4(n6263), .Q(round_key[100]));
   AO22X1 U7006 (.IN1(\key_mem[11][101] ), .IN2(n6491), .IN3(\key_mem[6][101] ), .IN4(
          n6476), .Q(n6267));
   AO221X1 U7007 (.IN1(\key_mem[4][101] ), .IN2(n6521), .IN3(\key_mem[5][101] ), .IN4(
          n6506), .IN5(n6267), .Q(n6273));
   AO222X1 U7008 (.IN1(\key_mem[9][101] ), .IN2(n6566), .IN3(\key_mem[8][101] ), .IN4(
          n6551), .IN5(\key_mem[10][101] ), .IN6(n6536), .Q(n6272));
   AO22X1 U7009 (.IN1(\key_mem[3][101] ), .IN2(n6596), .IN3(\key_mem[14][101] ), .IN4(
          n6581), .Q(n6268));
   AO221X1 U7010 (.IN1(\key_mem[12][101] ), .IN2(n6626), .IN3(\key_mem[13][101] ), .IN4(
          n6611), .IN5(n6268), .Q(n6271));
   AO22X1 U7011 (.IN1(\key_mem[7][101] ), .IN2(n6656), .IN3(\key_mem[2][101] ), .IN4(n6641)
          , .Q(n6269));
   AO221X1 U7012 (.IN1(\key_mem[0][101] ), .IN2(n6686), .IN3(\key_mem[1][101] ), .IN4(
          n6671), .IN5(n6269), .Q(n6270));
   OR4X1 U7013 (.IN1(n6273), .IN2(n6272), .IN3(n6271), .IN4(n6270), .Q(round_key[101]));
   AO22X1 U7014 (.IN1(\key_mem[11][102] ), .IN2(n6491), .IN3(\key_mem[6][102] ), .IN4(
          n6476), .Q(n6274));
   AO221X1 U7015 (.IN1(\key_mem[4][102] ), .IN2(n6521), .IN3(\key_mem[5][102] ), .IN4(
          n6506), .IN5(n6274), .Q(n6280));
   AO222X1 U7016 (.IN1(\key_mem[9][102] ), .IN2(n6566), .IN3(\key_mem[8][102] ), .IN4(
          n6551), .IN5(\key_mem[10][102] ), .IN6(n6536), .Q(n6279));
   AO22X1 U7017 (.IN1(\key_mem[3][102] ), .IN2(n6596), .IN3(\key_mem[14][102] ), .IN4(
          n6581), .Q(n6275));
   AO221X1 U7018 (.IN1(\key_mem[12][102] ), .IN2(n6626), .IN3(\key_mem[13][102] ), .IN4(
          n6611), .IN5(n6275), .Q(n6278));
   AO22X1 U7019 (.IN1(\key_mem[7][102] ), .IN2(n6656), .IN3(\key_mem[2][102] ), .IN4(n6641)
          , .Q(n6276));
   AO221X1 U7020 (.IN1(\key_mem[0][102] ), .IN2(n6686), .IN3(\key_mem[1][102] ), .IN4(
          n6671), .IN5(n6276), .Q(n6277));
   OR4X1 U7021 (.IN1(n6280), .IN2(n6279), .IN3(n6278), .IN4(n6277), .Q(round_key[102]));
   AO22X1 U7022 (.IN1(\key_mem[11][103] ), .IN2(n6491), .IN3(\key_mem[6][103] ), .IN4(
          n6476), .Q(n6281));
   AO221X1 U7023 (.IN1(\key_mem[4][103] ), .IN2(n6521), .IN3(\key_mem[5][103] ), .IN4(
          n6506), .IN5(n6281), .Q(n6287));
   AO222X1 U7024 (.IN1(\key_mem[9][103] ), .IN2(n6566), .IN3(\key_mem[8][103] ), .IN4(
          n6551), .IN5(\key_mem[10][103] ), .IN6(n6536), .Q(n6286));
   AO22X1 U7025 (.IN1(\key_mem[3][103] ), .IN2(n6596), .IN3(\key_mem[14][103] ), .IN4(
          n6581), .Q(n6282));
   AO221X1 U7026 (.IN1(\key_mem[12][103] ), .IN2(n6626), .IN3(\key_mem[13][103] ), .IN4(
          n6611), .IN5(n6282), .Q(n6285));
   AO22X1 U7027 (.IN1(\key_mem[7][103] ), .IN2(n6656), .IN3(\key_mem[2][103] ), .IN4(n6641)
          , .Q(n6283));
   AO221X1 U7028 (.IN1(\key_mem[0][103] ), .IN2(n6686), .IN3(\key_mem[1][103] ), .IN4(
          n6671), .IN5(n6283), .Q(n6284));
   OR4X1 U7029 (.IN1(n6287), .IN2(n6286), .IN3(n6285), .IN4(n6284), .Q(round_key[103]));
   AO22X1 U7030 (.IN1(\key_mem[11][104] ), .IN2(n6491), .IN3(\key_mem[6][104] ), .IN4(
          n6476), .Q(n6288));
   AO221X1 U7031 (.IN1(\key_mem[4][104] ), .IN2(n6521), .IN3(\key_mem[5][104] ), .IN4(
          n6506), .IN5(n6288), .Q(n6294));
   AO222X1 U7032 (.IN1(\key_mem[9][104] ), .IN2(n6566), .IN3(\key_mem[8][104] ), .IN4(
          n6551), .IN5(\key_mem[10][104] ), .IN6(n6536), .Q(n6293));
   AO22X1 U7033 (.IN1(\key_mem[3][104] ), .IN2(n6596), .IN3(\key_mem[14][104] ), .IN4(
          n6581), .Q(n6289));
   AO221X1 U7034 (.IN1(\key_mem[12][104] ), .IN2(n6626), .IN3(\key_mem[13][104] ), .IN4(
          n6611), .IN5(n6289), .Q(n6292));
   AO22X1 U7035 (.IN1(\key_mem[7][104] ), .IN2(n6656), .IN3(\key_mem[2][104] ), .IN4(n6641)
          , .Q(n6290));
   AO221X1 U7036 (.IN1(\key_mem[0][104] ), .IN2(n6686), .IN3(\key_mem[1][104] ), .IN4(
          n6671), .IN5(n6290), .Q(n6291));
   OR4X1 U7037 (.IN1(n6294), .IN2(n6293), .IN3(n6292), .IN4(n6291), .Q(round_key[104]));
   AO22X1 U7038 (.IN1(\key_mem[11][105] ), .IN2(n6491), .IN3(\key_mem[6][105] ), .IN4(
          n6476), .Q(n6295));
   AO221X1 U7039 (.IN1(\key_mem[4][105] ), .IN2(n6521), .IN3(\key_mem[5][105] ), .IN4(
          n6506), .IN5(n6295), .Q(n6301));
   AO222X1 U7040 (.IN1(\key_mem[9][105] ), .IN2(n6566), .IN3(\key_mem[8][105] ), .IN4(
          n6551), .IN5(\key_mem[10][105] ), .IN6(n6536), .Q(n6300));
   AO22X1 U7041 (.IN1(\key_mem[3][105] ), .IN2(n6596), .IN3(\key_mem[14][105] ), .IN4(
          n6581), .Q(n6296));
   AO221X1 U7042 (.IN1(\key_mem[12][105] ), .IN2(n6626), .IN3(\key_mem[13][105] ), .IN4(
          n6611), .IN5(n6296), .Q(n6299));
   AO22X1 U7043 (.IN1(\key_mem[7][105] ), .IN2(n6656), .IN3(\key_mem[2][105] ), .IN4(n6641)
          , .Q(n6297));
   AO221X1 U7044 (.IN1(\key_mem[0][105] ), .IN2(n6686), .IN3(\key_mem[1][105] ), .IN4(
          n6671), .IN5(n6297), .Q(n6298));
   OR4X1 U7045 (.IN1(n6301), .IN2(n6300), .IN3(n6299), .IN4(n6298), .Q(round_key[105]));
   AO22X1 U7046 (.IN1(\key_mem[11][106] ), .IN2(n6491), .IN3(\key_mem[6][106] ), .IN4(
          n6476), .Q(n6302));
   AO221X1 U7047 (.IN1(\key_mem[4][106] ), .IN2(n6521), .IN3(\key_mem[5][106] ), .IN4(
          n6506), .IN5(n6302), .Q(n6308));
   AO222X1 U7048 (.IN1(\key_mem[9][106] ), .IN2(n6566), .IN3(\key_mem[8][106] ), .IN4(
          n6551), .IN5(\key_mem[10][106] ), .IN6(n6536), .Q(n6307));
   AO22X1 U7049 (.IN1(\key_mem[3][106] ), .IN2(n6596), .IN3(\key_mem[14][106] ), .IN4(
          n6581), .Q(n6303));
   AO221X1 U7050 (.IN1(\key_mem[12][106] ), .IN2(n6626), .IN3(\key_mem[13][106] ), .IN4(
          n6611), .IN5(n6303), .Q(n6306));
   AO22X1 U7051 (.IN1(\key_mem[7][106] ), .IN2(n6656), .IN3(\key_mem[2][106] ), .IN4(n6641)
          , .Q(n6304));
   AO221X1 U7052 (.IN1(\key_mem[0][106] ), .IN2(n6686), .IN3(\key_mem[1][106] ), .IN4(
          n6671), .IN5(n6304), .Q(n6305));
   OR4X1 U7053 (.IN1(n6308), .IN2(n6307), .IN3(n6306), .IN4(n6305), .Q(round_key[106]));
   AO22X1 U7054 (.IN1(\key_mem[11][107] ), .IN2(n6491), .IN3(\key_mem[6][107] ), .IN4(
          n6476), .Q(n6309));
   AO221X1 U7055 (.IN1(\key_mem[4][107] ), .IN2(n6521), .IN3(\key_mem[5][107] ), .IN4(
          n6506), .IN5(n6309), .Q(n6315));
   AO222X1 U7056 (.IN1(\key_mem[9][107] ), .IN2(n6566), .IN3(\key_mem[8][107] ), .IN4(
          n6551), .IN5(\key_mem[10][107] ), .IN6(n6536), .Q(n6314));
   AO22X1 U7057 (.IN1(\key_mem[3][107] ), .IN2(n6596), .IN3(\key_mem[14][107] ), .IN4(
          n6581), .Q(n6310));
   AO221X1 U7058 (.IN1(\key_mem[12][107] ), .IN2(n6626), .IN3(\key_mem[13][107] ), .IN4(
          n6611), .IN5(n6310), .Q(n6313));
   AO22X1 U7059 (.IN1(\key_mem[7][107] ), .IN2(n6656), .IN3(\key_mem[2][107] ), .IN4(n6641)
          , .Q(n6311));
   AO221X1 U7060 (.IN1(\key_mem[0][107] ), .IN2(n6686), .IN3(\key_mem[1][107] ), .IN4(
          n6671), .IN5(n6311), .Q(n6312));
   OR4X1 U7061 (.IN1(n6315), .IN2(n6314), .IN3(n6313), .IN4(n6312), .Q(round_key[107]));
   AO22X1 U7062 (.IN1(\key_mem[11][108] ), .IN2(n6490), .IN3(\key_mem[6][108] ), .IN4(
          n6475), .Q(n6316));
   AO221X1 U7063 (.IN1(\key_mem[4][108] ), .IN2(n6520), .IN3(\key_mem[5][108] ), .IN4(
          n6505), .IN5(n6316), .Q(n6322));
   AO222X1 U7064 (.IN1(\key_mem[9][108] ), .IN2(n6565), .IN3(\key_mem[8][108] ), .IN4(
          n6550), .IN5(\key_mem[10][108] ), .IN6(n6535), .Q(n6321));
   AO22X1 U7065 (.IN1(\key_mem[3][108] ), .IN2(n6595), .IN3(\key_mem[14][108] ), .IN4(
          n6580), .Q(n6317));
   AO221X1 U7066 (.IN1(\key_mem[12][108] ), .IN2(n6625), .IN3(\key_mem[13][108] ), .IN4(
          n6610), .IN5(n6317), .Q(n6320));
   AO22X1 U7067 (.IN1(\key_mem[7][108] ), .IN2(n6655), .IN3(\key_mem[2][108] ), .IN4(n6640)
          , .Q(n6318));
   AO221X1 U7068 (.IN1(\key_mem[0][108] ), .IN2(n6685), .IN3(\key_mem[1][108] ), .IN4(
          n6670), .IN5(n6318), .Q(n6319));
   OR4X1 U7069 (.IN1(n6322), .IN2(n6321), .IN3(n6320), .IN4(n6319), .Q(round_key[108]));
   AO22X1 U7070 (.IN1(\key_mem[11][109] ), .IN2(n6490), .IN3(\key_mem[6][109] ), .IN4(
          n6475), .Q(n6323));
   AO221X1 U7071 (.IN1(\key_mem[4][109] ), .IN2(n6520), .IN3(\key_mem[5][109] ), .IN4(
          n6505), .IN5(n6323), .Q(n6329));
   AO222X1 U7072 (.IN1(\key_mem[9][109] ), .IN2(n6565), .IN3(\key_mem[8][109] ), .IN4(
          n6550), .IN5(\key_mem[10][109] ), .IN6(n6535), .Q(n6328));
   AO22X1 U7073 (.IN1(\key_mem[3][109] ), .IN2(n6595), .IN3(\key_mem[14][109] ), .IN4(
          n6580), .Q(n6324));
   AO221X1 U7074 (.IN1(\key_mem[12][109] ), .IN2(n6625), .IN3(\key_mem[13][109] ), .IN4(
          n6610), .IN5(n6324), .Q(n6327));
   AO22X1 U7075 (.IN1(\key_mem[7][109] ), .IN2(n6655), .IN3(\key_mem[2][109] ), .IN4(n6640)
          , .Q(n6325));
   AO221X1 U7076 (.IN1(\key_mem[0][109] ), .IN2(n6685), .IN3(\key_mem[1][109] ), .IN4(
          n6670), .IN5(n6325), .Q(n6326));
   OR4X1 U7077 (.IN1(n6329), .IN2(n6328), .IN3(n6327), .IN4(n6326), .Q(round_key[109]));
   AO22X1 U7078 (.IN1(\key_mem[11][110] ), .IN2(n6490), .IN3(\key_mem[6][110] ), .IN4(
          n6475), .Q(n6330));
   AO221X1 U7079 (.IN1(\key_mem[4][110] ), .IN2(n6520), .IN3(\key_mem[5][110] ), .IN4(
          n6505), .IN5(n6330), .Q(n6336));
   AO222X1 U7080 (.IN1(\key_mem[9][110] ), .IN2(n6565), .IN3(\key_mem[8][110] ), .IN4(
          n6550), .IN5(\key_mem[10][110] ), .IN6(n6535), .Q(n6335));
   AO22X1 U7081 (.IN1(\key_mem[3][110] ), .IN2(n6595), .IN3(\key_mem[14][110] ), .IN4(
          n6580), .Q(n6331));
   AO221X1 U7082 (.IN1(\key_mem[12][110] ), .IN2(n6625), .IN3(\key_mem[13][110] ), .IN4(
          n6610), .IN5(n6331), .Q(n6334));
   AO22X1 U7083 (.IN1(\key_mem[7][110] ), .IN2(n6655), .IN3(\key_mem[2][110] ), .IN4(n6640)
          , .Q(n6332));
   AO221X1 U7084 (.IN1(\key_mem[0][110] ), .IN2(n6685), .IN3(\key_mem[1][110] ), .IN4(
          n6670), .IN5(n6332), .Q(n6333));
   OR4X1 U7085 (.IN1(n6336), .IN2(n6335), .IN3(n6334), .IN4(n6333), .Q(round_key[110]));
   AO22X1 U7086 (.IN1(\key_mem[11][111] ), .IN2(n6490), .IN3(\key_mem[6][111] ), .IN4(
          n6475), .Q(n6337));
   AO221X1 U7087 (.IN1(\key_mem[4][111] ), .IN2(n6520), .IN3(\key_mem[5][111] ), .IN4(
          n6505), .IN5(n6337), .Q(n6343));
   AO222X1 U7088 (.IN1(\key_mem[9][111] ), .IN2(n6565), .IN3(\key_mem[8][111] ), .IN4(
          n6550), .IN5(\key_mem[10][111] ), .IN6(n6535), .Q(n6342));
   AO22X1 U7089 (.IN1(\key_mem[3][111] ), .IN2(n6595), .IN3(\key_mem[14][111] ), .IN4(
          n6580), .Q(n6338));
   AO221X1 U7090 (.IN1(\key_mem[12][111] ), .IN2(n6625), .IN3(\key_mem[13][111] ), .IN4(
          n6610), .IN5(n6338), .Q(n6341));
   AO22X1 U7091 (.IN1(\key_mem[7][111] ), .IN2(n6655), .IN3(\key_mem[2][111] ), .IN4(n6640)
          , .Q(n6339));
   AO221X1 U7092 (.IN1(\key_mem[0][111] ), .IN2(n6685), .IN3(\key_mem[1][111] ), .IN4(
          n6670), .IN5(n6339), .Q(n6340));
   OR4X1 U7093 (.IN1(n6343), .IN2(n6342), .IN3(n6341), .IN4(n6340), .Q(round_key[111]));
   AO22X1 U7094 (.IN1(\key_mem[11][112] ), .IN2(n6490), .IN3(\key_mem[6][112] ), .IN4(
          n6475), .Q(n6344));
   AO221X1 U7095 (.IN1(\key_mem[4][112] ), .IN2(n6520), .IN3(\key_mem[5][112] ), .IN4(
          n6505), .IN5(n6344), .Q(n6350));
   AO222X1 U7096 (.IN1(\key_mem[9][112] ), .IN2(n6565), .IN3(\key_mem[8][112] ), .IN4(
          n6550), .IN5(\key_mem[10][112] ), .IN6(n6535), .Q(n6349));
   AO22X1 U7097 (.IN1(\key_mem[3][112] ), .IN2(n6595), .IN3(\key_mem[14][112] ), .IN4(
          n6580), .Q(n6345));
   AO221X1 U7098 (.IN1(\key_mem[12][112] ), .IN2(n6625), .IN3(\key_mem[13][112] ), .IN4(
          n6610), .IN5(n6345), .Q(n6348));
   AO22X1 U7099 (.IN1(\key_mem[7][112] ), .IN2(n6655), .IN3(\key_mem[2][112] ), .IN4(n6640)
          , .Q(n6346));
   AO221X1 U7100 (.IN1(\key_mem[0][112] ), .IN2(n6685), .IN3(\key_mem[1][112] ), .IN4(
          n6670), .IN5(n6346), .Q(n6347));
   OR4X1 U7101 (.IN1(n6350), .IN2(n6349), .IN3(n6348), .IN4(n6347), .Q(round_key[112]));
   AO22X1 U7102 (.IN1(\key_mem[11][113] ), .IN2(n6490), .IN3(\key_mem[6][113] ), .IN4(
          n6475), .Q(n6351));
   AO221X1 U7103 (.IN1(\key_mem[4][113] ), .IN2(n6520), .IN3(\key_mem[5][113] ), .IN4(
          n6505), .IN5(n6351), .Q(n6357));
   AO222X1 U7104 (.IN1(\key_mem[9][113] ), .IN2(n6565), .IN3(\key_mem[8][113] ), .IN4(
          n6550), .IN5(\key_mem[10][113] ), .IN6(n6535), .Q(n6356));
   AO22X1 U7105 (.IN1(\key_mem[3][113] ), .IN2(n6595), .IN3(\key_mem[14][113] ), .IN4(
          n6580), .Q(n6352));
   AO221X1 U7106 (.IN1(\key_mem[12][113] ), .IN2(n6625), .IN3(\key_mem[13][113] ), .IN4(
          n6610), .IN5(n6352), .Q(n6355));
   AO22X1 U7107 (.IN1(\key_mem[7][113] ), .IN2(n6655), .IN3(\key_mem[2][113] ), .IN4(n6640)
          , .Q(n6353));
   AO221X1 U7108 (.IN1(\key_mem[0][113] ), .IN2(n6685), .IN3(\key_mem[1][113] ), .IN4(
          n6670), .IN5(n6353), .Q(n6354));
   OR4X1 U7109 (.IN1(n6357), .IN2(n6356), .IN3(n6355), .IN4(n6354), .Q(round_key[113]));
   AO22X1 U7110 (.IN1(\key_mem[11][114] ), .IN2(n6490), .IN3(\key_mem[6][114] ), .IN4(
          n6475), .Q(n6358));
   AO221X1 U7111 (.IN1(\key_mem[4][114] ), .IN2(n6520), .IN3(\key_mem[5][114] ), .IN4(
          n6505), .IN5(n6358), .Q(n6364));
   AO222X1 U7112 (.IN1(\key_mem[9][114] ), .IN2(n6565), .IN3(\key_mem[8][114] ), .IN4(
          n6550), .IN5(\key_mem[10][114] ), .IN6(n6535), .Q(n6363));
   AO22X1 U7113 (.IN1(\key_mem[3][114] ), .IN2(n6595), .IN3(\key_mem[14][114] ), .IN4(
          n6580), .Q(n6359));
   AO221X1 U7114 (.IN1(\key_mem[12][114] ), .IN2(n6625), .IN3(\key_mem[13][114] ), .IN4(
          n6610), .IN5(n6359), .Q(n6362));
   AO22X1 U7115 (.IN1(\key_mem[7][114] ), .IN2(n6655), .IN3(\key_mem[2][114] ), .IN4(n6640)
          , .Q(n6360));
   AO221X1 U7116 (.IN1(\key_mem[0][114] ), .IN2(n6685), .IN3(\key_mem[1][114] ), .IN4(
          n6670), .IN5(n6360), .Q(n6361));
   OR4X1 U7117 (.IN1(n6364), .IN2(n6363), .IN3(n6362), .IN4(n6361), .Q(round_key[114]));
   AO22X1 U7118 (.IN1(\key_mem[11][115] ), .IN2(n6490), .IN3(\key_mem[6][115] ), .IN4(
          n6475), .Q(n6365));
   AO221X1 U7119 (.IN1(\key_mem[4][115] ), .IN2(n6520), .IN3(\key_mem[5][115] ), .IN4(
          n6505), .IN5(n6365), .Q(n6371));
   AO222X1 U7120 (.IN1(\key_mem[9][115] ), .IN2(n6565), .IN3(\key_mem[8][115] ), .IN4(
          n6550), .IN5(\key_mem[10][115] ), .IN6(n6535), .Q(n6370));
   AO22X1 U7121 (.IN1(\key_mem[3][115] ), .IN2(n6595), .IN3(\key_mem[14][115] ), .IN4(
          n6580), .Q(n6366));
   AO221X1 U7122 (.IN1(\key_mem[12][115] ), .IN2(n6625), .IN3(\key_mem[13][115] ), .IN4(
          n6610), .IN5(n6366), .Q(n6369));
   AO22X1 U7123 (.IN1(\key_mem[7][115] ), .IN2(n6655), .IN3(\key_mem[2][115] ), .IN4(n6640)
          , .Q(n6367));
   AO221X1 U7124 (.IN1(\key_mem[0][115] ), .IN2(n6685), .IN3(\key_mem[1][115] ), .IN4(
          n6670), .IN5(n6367), .Q(n6368));
   OR4X1 U7125 (.IN1(n6371), .IN2(n6370), .IN3(n6369), .IN4(n6368), .Q(round_key[115]));
   AO22X1 U7126 (.IN1(\key_mem[11][116] ), .IN2(n6490), .IN3(\key_mem[6][116] ), .IN4(
          n6475), .Q(n6372));
   AO221X1 U7127 (.IN1(\key_mem[4][116] ), .IN2(n6520), .IN3(\key_mem[5][116] ), .IN4(
          n6505), .IN5(n6372), .Q(n6378));
   AO222X1 U7128 (.IN1(\key_mem[9][116] ), .IN2(n6565), .IN3(\key_mem[8][116] ), .IN4(
          n6550), .IN5(\key_mem[10][116] ), .IN6(n6535), .Q(n6377));
   AO22X1 U7129 (.IN1(\key_mem[3][116] ), .IN2(n6595), .IN3(\key_mem[14][116] ), .IN4(
          n6580), .Q(n6373));
   AO221X1 U7130 (.IN1(\key_mem[12][116] ), .IN2(n6625), .IN3(\key_mem[13][116] ), .IN4(
          n6610), .IN5(n6373), .Q(n6376));
   AO22X1 U7131 (.IN1(\key_mem[7][116] ), .IN2(n6655), .IN3(\key_mem[2][116] ), .IN4(n6640)
          , .Q(n6374));
   AO221X1 U7132 (.IN1(\key_mem[0][116] ), .IN2(n6685), .IN3(\key_mem[1][116] ), .IN4(
          n6670), .IN5(n6374), .Q(n6375));
   OR4X1 U7133 (.IN1(n6378), .IN2(n6377), .IN3(n6376), .IN4(n6375), .Q(round_key[116]));
   AO22X1 U7134 (.IN1(\key_mem[11][117] ), .IN2(n6490), .IN3(\key_mem[6][117] ), .IN4(
          n6475), .Q(n6379));
   AO221X1 U7135 (.IN1(\key_mem[4][117] ), .IN2(n6520), .IN3(\key_mem[5][117] ), .IN4(
          n6505), .IN5(n6379), .Q(n6385));
   AO222X1 U7136 (.IN1(\key_mem[9][117] ), .IN2(n6565), .IN3(\key_mem[8][117] ), .IN4(
          n6550), .IN5(\key_mem[10][117] ), .IN6(n6535), .Q(n6384));
   AO22X1 U7137 (.IN1(\key_mem[3][117] ), .IN2(n6595), .IN3(\key_mem[14][117] ), .IN4(
          n6580), .Q(n6380));
   AO221X1 U7138 (.IN1(\key_mem[12][117] ), .IN2(n6625), .IN3(\key_mem[13][117] ), .IN4(
          n6610), .IN5(n6380), .Q(n6383));
   AO22X1 U7139 (.IN1(\key_mem[7][117] ), .IN2(n6655), .IN3(\key_mem[2][117] ), .IN4(n6640)
          , .Q(n6381));
   AO221X1 U7140 (.IN1(\key_mem[0][117] ), .IN2(n6685), .IN3(\key_mem[1][117] ), .IN4(
          n6670), .IN5(n6381), .Q(n6382));
   OR4X1 U7141 (.IN1(n6385), .IN2(n6384), .IN3(n6383), .IN4(n6382), .Q(round_key[117]));
   AO22X1 U7142 (.IN1(\key_mem[11][118] ), .IN2(n6490), .IN3(\key_mem[6][118] ), .IN4(
          n6475), .Q(n6386));
   AO221X1 U7143 (.IN1(\key_mem[4][118] ), .IN2(n6520), .IN3(\key_mem[5][118] ), .IN4(
          n6505), .IN5(n6386), .Q(n6392));
   AO222X1 U7144 (.IN1(\key_mem[9][118] ), .IN2(n6565), .IN3(\key_mem[8][118] ), .IN4(
          n6550), .IN5(\key_mem[10][118] ), .IN6(n6535), .Q(n6391));
   AO22X1 U7145 (.IN1(\key_mem[3][118] ), .IN2(n6595), .IN3(\key_mem[14][118] ), .IN4(
          n6580), .Q(n6387));
   AO221X1 U7146 (.IN1(\key_mem[12][118] ), .IN2(n6625), .IN3(\key_mem[13][118] ), .IN4(
          n6610), .IN5(n6387), .Q(n6390));
   AO22X1 U7147 (.IN1(\key_mem[7][118] ), .IN2(n6655), .IN3(\key_mem[2][118] ), .IN4(n6640)
          , .Q(n6388));
   AO221X1 U7148 (.IN1(\key_mem[0][118] ), .IN2(n6685), .IN3(\key_mem[1][118] ), .IN4(
          n6670), .IN5(n6388), .Q(n6389));
   OR4X1 U7149 (.IN1(n6392), .IN2(n6391), .IN3(n6390), .IN4(n6389), .Q(round_key[118]));
   AO22X1 U7150 (.IN1(\key_mem[11][119] ), .IN2(n6490), .IN3(\key_mem[6][119] ), .IN4(
          n6475), .Q(n6393));
   AO221X1 U7151 (.IN1(\key_mem[4][119] ), .IN2(n6520), .IN3(\key_mem[5][119] ), .IN4(
          n6505), .IN5(n6393), .Q(n6399));
   AO222X1 U7152 (.IN1(\key_mem[9][119] ), .IN2(n6565), .IN3(\key_mem[8][119] ), .IN4(
          n6550), .IN5(\key_mem[10][119] ), .IN6(n6535), .Q(n6398));
   AO22X1 U7153 (.IN1(\key_mem[3][119] ), .IN2(n6595), .IN3(\key_mem[14][119] ), .IN4(
          n6580), .Q(n6394));
   AO221X1 U7154 (.IN1(\key_mem[12][119] ), .IN2(n6625), .IN3(\key_mem[13][119] ), .IN4(
          n6610), .IN5(n6394), .Q(n6397));
   AO22X1 U7155 (.IN1(\key_mem[7][119] ), .IN2(n6655), .IN3(\key_mem[2][119] ), .IN4(n6640)
          , .Q(n6395));
   AO221X1 U7156 (.IN1(\key_mem[0][119] ), .IN2(n6685), .IN3(\key_mem[1][119] ), .IN4(
          n6670), .IN5(n6395), .Q(n6396));
   OR4X1 U7157 (.IN1(n6399), .IN2(n6398), .IN3(n6397), .IN4(n6396), .Q(round_key[119]));
   AO22X1 U7158 (.IN1(\key_mem[11][120] ), .IN2(n6489), .IN3(\key_mem[6][120] ), .IN4(
          n6474), .Q(n6400));
   AO221X1 U7159 (.IN1(\key_mem[4][120] ), .IN2(n6519), .IN3(\key_mem[5][120] ), .IN4(
          n6504), .IN5(n6400), .Q(n6406));
   AO222X1 U7160 (.IN1(\key_mem[9][120] ), .IN2(n6564), .IN3(\key_mem[8][120] ), .IN4(
          n6549), .IN5(\key_mem[10][120] ), .IN6(n6534), .Q(n6405));
   AO22X1 U7161 (.IN1(\key_mem[3][120] ), .IN2(n6594), .IN3(\key_mem[14][120] ), .IN4(
          n6579), .Q(n6401));
   AO221X1 U7162 (.IN1(\key_mem[12][120] ), .IN2(n6624), .IN3(\key_mem[13][120] ), .IN4(
          n6609), .IN5(n6401), .Q(n6404));
   AO22X1 U7163 (.IN1(\key_mem[7][120] ), .IN2(n6654), .IN3(\key_mem[2][120] ), .IN4(n6639)
          , .Q(n6402));
   AO221X1 U7164 (.IN1(\key_mem[0][120] ), .IN2(n6684), .IN3(\key_mem[1][120] ), .IN4(
          n6669), .IN5(n6402), .Q(n6403));
   OR4X1 U7165 (.IN1(n6406), .IN2(n6405), .IN3(n6404), .IN4(n6403), .Q(round_key[120]));
   AO22X1 U7166 (.IN1(\key_mem[11][121] ), .IN2(n6489), .IN3(\key_mem[6][121] ), .IN4(
          n6474), .Q(n6407));
   AO221X1 U7167 (.IN1(\key_mem[4][121] ), .IN2(n6519), .IN3(\key_mem[5][121] ), .IN4(
          n6504), .IN5(n6407), .Q(n6413));
   AO222X1 U7168 (.IN1(\key_mem[9][121] ), .IN2(n6564), .IN3(\key_mem[8][121] ), .IN4(
          n6549), .IN5(\key_mem[10][121] ), .IN6(n6534), .Q(n6412));
   AO22X1 U7169 (.IN1(\key_mem[3][121] ), .IN2(n6594), .IN3(\key_mem[14][121] ), .IN4(
          n6579), .Q(n6408));
   AO221X1 U7170 (.IN1(\key_mem[12][121] ), .IN2(n6624), .IN3(\key_mem[13][121] ), .IN4(
          n6609), .IN5(n6408), .Q(n6411));
   AO22X1 U7171 (.IN1(\key_mem[7][121] ), .IN2(n6654), .IN3(\key_mem[2][121] ), .IN4(n6639)
          , .Q(n6409));
   AO221X1 U7172 (.IN1(\key_mem[0][121] ), .IN2(n6684), .IN3(\key_mem[1][121] ), .IN4(
          n6669), .IN5(n6409), .Q(n6410));
   OR4X1 U7173 (.IN1(n6413), .IN2(n6412), .IN3(n6411), .IN4(n6410), .Q(round_key[121]));
   AO22X1 U7174 (.IN1(\key_mem[11][122] ), .IN2(n6489), .IN3(\key_mem[6][122] ), .IN4(
          n6474), .Q(n6414));
   AO221X1 U7175 (.IN1(\key_mem[4][122] ), .IN2(n6519), .IN3(\key_mem[5][122] ), .IN4(
          n6504), .IN5(n6414), .Q(n6420));
   AO222X1 U7176 (.IN1(\key_mem[9][122] ), .IN2(n6564), .IN3(\key_mem[8][122] ), .IN4(
          n6549), .IN5(\key_mem[10][122] ), .IN6(n6534), .Q(n6419));
   AO22X1 U7177 (.IN1(\key_mem[3][122] ), .IN2(n6594), .IN3(\key_mem[14][122] ), .IN4(
          n6579), .Q(n6415));
   AO221X1 U7178 (.IN1(\key_mem[12][122] ), .IN2(n6624), .IN3(\key_mem[13][122] ), .IN4(
          n6609), .IN5(n6415), .Q(n6418));
   AO22X1 U7179 (.IN1(\key_mem[7][122] ), .IN2(n6654), .IN3(\key_mem[2][122] ), .IN4(n6639)
          , .Q(n6416));
   AO221X1 U7180 (.IN1(\key_mem[0][122] ), .IN2(n6684), .IN3(\key_mem[1][122] ), .IN4(
          n6669), .IN5(n6416), .Q(n6417));
   OR4X1 U7181 (.IN1(n6420), .IN2(n6419), .IN3(n6418), .IN4(n6417), .Q(round_key[122]));
   AO22X1 U7182 (.IN1(\key_mem[11][123] ), .IN2(n6489), .IN3(\key_mem[6][123] ), .IN4(
          n6474), .Q(n6421));
   AO221X1 U7183 (.IN1(\key_mem[4][123] ), .IN2(n6519), .IN3(\key_mem[5][123] ), .IN4(
          n6504), .IN5(n6421), .Q(n6427));
   AO222X1 U7184 (.IN1(\key_mem[9][123] ), .IN2(n6564), .IN3(\key_mem[8][123] ), .IN4(
          n6549), .IN5(\key_mem[10][123] ), .IN6(n6534), .Q(n6426));
   AO22X1 U7185 (.IN1(\key_mem[3][123] ), .IN2(n6594), .IN3(\key_mem[14][123] ), .IN4(
          n6579), .Q(n6422));
   AO221X1 U7186 (.IN1(\key_mem[12][123] ), .IN2(n6624), .IN3(\key_mem[13][123] ), .IN4(
          n6609), .IN5(n6422), .Q(n6425));
   AO22X1 U7187 (.IN1(\key_mem[7][123] ), .IN2(n6654), .IN3(\key_mem[2][123] ), .IN4(n6639)
          , .Q(n6423));
   AO221X1 U7188 (.IN1(\key_mem[0][123] ), .IN2(n6684), .IN3(\key_mem[1][123] ), .IN4(
          n6669), .IN5(n6423), .Q(n6424));
   OR4X1 U7189 (.IN1(n6427), .IN2(n6426), .IN3(n6425), .IN4(n6424), .Q(round_key[123]));
   AO22X1 U7190 (.IN1(\key_mem[11][124] ), .IN2(n6489), .IN3(\key_mem[6][124] ), .IN4(
          n6474), .Q(n6428));
   AO221X1 U7191 (.IN1(\key_mem[4][124] ), .IN2(n6519), .IN3(\key_mem[5][124] ), .IN4(
          n6504), .IN5(n6428), .Q(n6434));
   AO222X1 U7192 (.IN1(\key_mem[9][124] ), .IN2(n6564), .IN3(\key_mem[8][124] ), .IN4(
          n6549), .IN5(\key_mem[10][124] ), .IN6(n6534), .Q(n6433));
   AO22X1 U7193 (.IN1(\key_mem[3][124] ), .IN2(n6594), .IN3(\key_mem[14][124] ), .IN4(
          n6579), .Q(n6429));
   AO221X1 U7194 (.IN1(\key_mem[12][124] ), .IN2(n6624), .IN3(\key_mem[13][124] ), .IN4(
          n6609), .IN5(n6429), .Q(n6432));
   AO22X1 U7195 (.IN1(\key_mem[7][124] ), .IN2(n6654), .IN3(\key_mem[2][124] ), .IN4(n6639)
          , .Q(n6430));
   AO221X1 U7196 (.IN1(\key_mem[0][124] ), .IN2(n6684), .IN3(\key_mem[1][124] ), .IN4(
          n6669), .IN5(n6430), .Q(n6431));
   OR4X1 U7197 (.IN1(n6434), .IN2(n6433), .IN3(n6432), .IN4(n6431), .Q(round_key[124]));
   AO22X1 U7198 (.IN1(\key_mem[11][125] ), .IN2(n6489), .IN3(\key_mem[6][125] ), .IN4(
          n6474), .Q(n6435));
   AO221X1 U7199 (.IN1(\key_mem[4][125] ), .IN2(n6519), .IN3(\key_mem[5][125] ), .IN4(
          n6504), .IN5(n6435), .Q(n6441));
   AO222X1 U7200 (.IN1(\key_mem[9][125] ), .IN2(n6564), .IN3(\key_mem[8][125] ), .IN4(
          n6549), .IN5(\key_mem[10][125] ), .IN6(n6534), .Q(n6440));
   AO22X1 U7201 (.IN1(\key_mem[3][125] ), .IN2(n6594), .IN3(\key_mem[14][125] ), .IN4(
          n6579), .Q(n6436));
   AO221X1 U7202 (.IN1(\key_mem[12][125] ), .IN2(n6624), .IN3(\key_mem[13][125] ), .IN4(
          n6609), .IN5(n6436), .Q(n6439));
   AO22X1 U7203 (.IN1(\key_mem[7][125] ), .IN2(n6654), .IN3(\key_mem[2][125] ), .IN4(n6639)
          , .Q(n6437));
   AO221X1 U7204 (.IN1(\key_mem[0][125] ), .IN2(n6684), .IN3(\key_mem[1][125] ), .IN4(
          n6669), .IN5(n6437), .Q(n6438));
   OR4X1 U7205 (.IN1(n6441), .IN2(n6440), .IN3(n6439), .IN4(n6438), .Q(round_key[125]));
   AO22X1 U7206 (.IN1(\key_mem[11][126] ), .IN2(n6489), .IN3(\key_mem[6][126] ), .IN4(
          n6474), .Q(n6442));
   AO221X1 U7207 (.IN1(\key_mem[4][126] ), .IN2(n6519), .IN3(\key_mem[5][126] ), .IN4(
          n6504), .IN5(n6442), .Q(n6448));
   AO222X1 U7208 (.IN1(\key_mem[9][126] ), .IN2(n6564), .IN3(\key_mem[8][126] ), .IN4(
          n6549), .IN5(\key_mem[10][126] ), .IN6(n6534), .Q(n6447));
   AO22X1 U7209 (.IN1(\key_mem[3][126] ), .IN2(n6594), .IN3(\key_mem[14][126] ), .IN4(
          n6579), .Q(n6443));
   AO221X1 U7210 (.IN1(\key_mem[12][126] ), .IN2(n6624), .IN3(\key_mem[13][126] ), .IN4(
          n6609), .IN5(n6443), .Q(n6446));
   AO22X1 U7211 (.IN1(\key_mem[7][126] ), .IN2(n6654), .IN3(\key_mem[2][126] ), .IN4(n6639)
          , .Q(n6444));
   AO221X1 U7212 (.IN1(\key_mem[0][126] ), .IN2(n6684), .IN3(\key_mem[1][126] ), .IN4(
          n6669), .IN5(n6444), .Q(n6445));
   OR4X1 U7213 (.IN1(n6448), .IN2(n6447), .IN3(n6446), .IN4(n6445), .Q(round_key[126]));
   AO22X1 U7214 (.IN1(\key_mem[11][127] ), .IN2(n6489), .IN3(\key_mem[6][127] ), .IN4(
          n6474), .Q(n6451));
   AO221X1 U7215 (.IN1(\key_mem[4][127] ), .IN2(n6519), .IN3(\key_mem[5][127] ), .IN4(
          n6504), .IN5(n6451), .Q(n6470));
   AO222X1 U7216 (.IN1(\key_mem[9][127] ), .IN2(n6564), .IN3(\key_mem[8][127] ), .IN4(
          n6549), .IN5(\key_mem[10][127] ), .IN6(n6534), .Q(n6469));
   AO22X1 U7217 (.IN1(\key_mem[3][127] ), .IN2(n6594), .IN3(\key_mem[14][127] ), .IN4(
          n6579), .Q(n6459));
   AO221X1 U7218 (.IN1(\key_mem[12][127] ), .IN2(n6624), .IN3(\key_mem[13][127] ), .IN4(
          n6609), .IN5(n6459), .Q(n6468));
   AO22X1 U7219 (.IN1(\key_mem[7][127] ), .IN2(n6654), .IN3(\key_mem[2][127] ), .IN4(n6639)
          , .Q(n6464));
   AO221X1 U7220 (.IN1(\key_mem[0][127] ), .IN2(n6684), .IN3(\key_mem[1][127] ), .IN4(
          n6669), .IN5(n6464), .Q(n6467));
   OR4X1 U7221 (.IN1(n6470), .IN2(n6469), .IN3(n6468), .IN4(n6467), .Q(round_key[127]));
   NBUFFX2 U7222 (.INP(n6462), .Z(n6652));
   NBUFFX2 U7223 (.INP(n6462), .Z(n6653));
   AND2X2 U7224 (.IN1(n2233), .IN2(n2232), .Q(n6462));
   AO22X1 U7225 (.IN1(n6813), .IN2(n2340), .IN3(\key_mem[1][118] ), .IN4(n6822), .Q(n3562)
          );
   INVX0 U7226 (.INP(n2945), .ZN(n6702));
   INVX0 U7227 (.INP(n6702), .ZN(n6703));
   INVX0 U7228 (.INP(n6702), .ZN(n6704));
   INVX0 U7229 (.INP(n6702), .ZN(n6705));
   INVX0 U7230 (.INP(n6702), .ZN(n6706));
   INVX0 U7231 (.INP(n6702), .ZN(n6707));
   INVX0 U7232 (.INP(n6702), .ZN(n6708));
   INVX0 U7233 (.INP(n6702), .ZN(n6709));
   INVX0 U7234 (.INP(n6702), .ZN(n6710));
   INVX0 U7235 (.INP(n6702), .ZN(n6711));
   INVX0 U7236 (.INP(n6830), .ZN(n6829));
   INVX0 U7237 (.INP(n6836), .ZN(n6835));
   INVX0 U7238 (.INP(n6841), .ZN(n6840));
   INVX0 U7239 (.INP(n6828), .ZN(n6827));
   INVX0 U7240 (.INP(n6828), .ZN(n6826));
   INVX0 U7241 (.INP(n6833), .ZN(n6832));
   INVX0 U7242 (.INP(n6834), .ZN(n6831));
   INVX0 U7243 (.INP(n6839), .ZN(n6837));
   INVX0 U7244 (.INP(n7186), .ZN(n6830));
   INVX0 U7245 (.INP(n6987), .ZN(n6841));
   INVX0 U7246 (.INP(n6986), .ZN(n6836));
   INVX0 U7247 (.INP(n6829), .ZN(n6828));
   INVX0 U7248 (.INP(n6835), .ZN(n6833));
   INVX0 U7249 (.INP(n6835), .ZN(n6834));
   INVX0 U7250 (.INP(n6840), .ZN(n6838));
   INVX0 U7251 (.INP(n6840), .ZN(n6839));
   AND3X1 U7252 (.IN1(n2931), .IN2(n2212), .IN3(n2934), .Q(n6990));
   INVX0 U7253 (.INP(n7284), .ZN(n6916));
   INVX0 U7254 (.INP(n7285), .ZN(n6920));
   INVX0 U7255 (.INP(n6925), .ZN(n6924));
   INVX0 U7256 (.INP(n7021), .ZN(n6886));
   INVX0 U7257 (.INP(n7021), .ZN(n6887));
   INVX0 U7258 (.INP(n6923), .ZN(n6922));
   INVX0 U7259 (.INP(n6923), .ZN(n6921));
   INVX0 U7260 (.INP(n7285), .ZN(n6888));
   INVX0 U7261 (.INP(n6925), .ZN(n6889));
   INVX0 U7262 (.INP(n6990), .ZN(n6925));
   INVX0 U7263 (.INP(n7022), .ZN(n6890));
   INVX0 U7264 (.INP(n6920), .ZN(n6919));
   INVX0 U7265 (.INP(n6916), .ZN(n6918));
   INVX0 U7266 (.INP(n6889), .ZN(n6914));
   INVX0 U7267 (.INP(n6916), .ZN(n6915));
   INVX0 U7268 (.INP(n6889), .ZN(n6917));
   INVX0 U7269 (.INP(n6924), .ZN(n6923));
   INVX0 U7270 (.INP(n7010), .ZN(n6712));
   INVX0 U7271 (.INP(n7228), .ZN(n6713));
   INVX0 U7272 (.INP(n6713), .ZN(n6714));
   INVX0 U7273 (.INP(n6713), .ZN(n6715));
   INVX0 U7274 (.INP(n6713), .ZN(n6716));
   INVX0 U7275 (.INP(n7230), .ZN(n6717));
   INVX0 U7276 (.INP(n6723), .ZN(n6718));
   INVX0 U7277 (.INP(n6748), .ZN(n6719));
   INVX0 U7278 (.INP(n6751), .ZN(n6720));
   INVX0 U7279 (.INP(n7230), .ZN(n6721));
   INVX0 U7280 (.INP(n6749), .ZN(n6722));
   INVX0 U7281 (.INP(n7229), .ZN(n6723));
   INVX0 U7282 (.INP(n6723), .ZN(n6724));
   INVX0 U7283 (.INP(n6723), .ZN(n6725));
   INVX0 U7284 (.INP(n6713), .ZN(n6726));
   INVX0 U7285 (.INP(n6723), .ZN(n6727));
   INVX0 U7286 (.INP(n6885), .ZN(n6728));
   INVX0 U7287 (.INP(n6728), .ZN(n6729));
   INVX0 U7288 (.INP(n6728), .ZN(n6730));
   INVX0 U7289 (.INP(n6728), .ZN(n6731));
   INVX0 U7290 (.INP(n6910), .ZN(n6732));
   INVX0 U7291 (.INP(n6732), .ZN(n6733));
   INVX0 U7292 (.INP(n6732), .ZN(n6734));
   INVX0 U7293 (.INP(n6732), .ZN(n6735));
   INVX0 U7294 (.INP(n6911), .ZN(n6736));
   INVX0 U7295 (.INP(n6736), .ZN(n6737));
   INVX0 U7296 (.INP(n6736), .ZN(n6738));
   INVX0 U7297 (.INP(n6736), .ZN(n6739));
   INVX0 U7298 (.INP(n6883), .ZN(n6740));
   INVX0 U7299 (.INP(n6740), .ZN(n6741));
   INVX0 U7300 (.INP(n6740), .ZN(n6742));
   INVX0 U7301 (.INP(n6740), .ZN(n6743));
   INVX0 U7302 (.INP(n6882), .ZN(n6744));
   INVX0 U7303 (.INP(n6744), .ZN(n6745));
   INVX0 U7304 (.INP(n6744), .ZN(n6746));
   INVX0 U7305 (.INP(n6744), .ZN(n6747));
   INVX0 U7306 (.INP(n7234), .ZN(n6748));
   INVX0 U7307 (.INP(n7234), .ZN(n6749));
   INVX0 U7308 (.INP(n7234), .ZN(n6750));
   INVX0 U7309 (.INP(n7234), .ZN(n6751));
   INVX0 U7310 (.INP(n7234), .ZN(n6752));
   INVX0 U7311 (.INP(n6712), .ZN(n6753));
   INVX0 U7312 (.INP(n6753), .ZN(n6754));
   INVX0 U7313 (.INP(n6753), .ZN(n6755));
   INVX0 U7314 (.INP(n6753), .ZN(n6756));
   INVX0 U7315 (.INP(n6753), .ZN(n6757));
   INVX0 U7316 (.INP(n6753), .ZN(n6758));
   INVX0 U7317 (.INP(n6913), .ZN(n6912));
   INVX0 U7318 (.INP(n6885), .ZN(n6884));
   INVX0 U7319 (.INP(n7232), .ZN(n6913));
   INVX0 U7320 (.INP(n7011), .ZN(n6885));
   INVX0 U7321 (.INP(n6912), .ZN(n6910));
   INVX0 U7322 (.INP(n6912), .ZN(n6911));
   INVX0 U7323 (.INP(n6884), .ZN(n6883));
   INVX0 U7324 (.INP(n6884), .ZN(n6882));
   INVX0 U7325 (.INP(n7005), .ZN(n6759));
   INVX0 U7326 (.INP(n7204), .ZN(n6760));
   INVX0 U7327 (.INP(n6760), .ZN(n6761));
   INVX0 U7328 (.INP(n6760), .ZN(n6762));
   INVX0 U7329 (.INP(n6760), .ZN(n6763));
   INVX0 U7330 (.INP(n7206), .ZN(n6764));
   INVX0 U7331 (.INP(n6770), .ZN(n6765));
   INVX0 U7332 (.INP(n6795), .ZN(n6766));
   INVX0 U7333 (.INP(n6798), .ZN(n6767));
   INVX0 U7334 (.INP(n7206), .ZN(n6768));
   INVX0 U7335 (.INP(n6796), .ZN(n6769));
   INVX0 U7336 (.INP(n7205), .ZN(n6770));
   INVX0 U7337 (.INP(n6770), .ZN(n6771));
   INVX0 U7338 (.INP(n6770), .ZN(n6772));
   INVX0 U7339 (.INP(n6760), .ZN(n6773));
   INVX0 U7340 (.INP(n6770), .ZN(n6774));
   INVX0 U7341 (.INP(n6881), .ZN(n6775));
   INVX0 U7342 (.INP(n6775), .ZN(n6776));
   INVX0 U7343 (.INP(n6775), .ZN(n6777));
   INVX0 U7344 (.INP(n6775), .ZN(n6778));
   INVX0 U7345 (.INP(n6906), .ZN(n6779));
   INVX0 U7346 (.INP(n6779), .ZN(n6780));
   INVX0 U7347 (.INP(n6779), .ZN(n6781));
   INVX0 U7348 (.INP(n6779), .ZN(n6782));
   INVX0 U7349 (.INP(n6907), .ZN(n6783));
   INVX0 U7350 (.INP(n6783), .ZN(n6784));
   INVX0 U7351 (.INP(n6783), .ZN(n6785));
   INVX0 U7352 (.INP(n6783), .ZN(n6786));
   INVX0 U7353 (.INP(n6879), .ZN(n6787));
   INVX0 U7354 (.INP(n6787), .ZN(n6788));
   INVX0 U7355 (.INP(n6787), .ZN(n6789));
   INVX0 U7356 (.INP(n6787), .ZN(n6790));
   INVX0 U7357 (.INP(n6878), .ZN(n6791));
   INVX0 U7358 (.INP(n6791), .ZN(n6792));
   INVX0 U7359 (.INP(n6791), .ZN(n6793));
   INVX0 U7360 (.INP(n6791), .ZN(n6794));
   INVX0 U7361 (.INP(n7210), .ZN(n6795));
   INVX0 U7362 (.INP(n7210), .ZN(n6796));
   INVX0 U7363 (.INP(n7210), .ZN(n6797));
   INVX0 U7364 (.INP(n7210), .ZN(n6798));
   INVX0 U7365 (.INP(n7210), .ZN(n6799));
   INVX0 U7366 (.INP(n6759), .ZN(n6800));
   INVX0 U7367 (.INP(n6800), .ZN(n6801));
   INVX0 U7368 (.INP(n6800), .ZN(n6802));
   INVX0 U7369 (.INP(n6800), .ZN(n6803));
   INVX0 U7370 (.INP(n6800), .ZN(n6804));
   INVX0 U7371 (.INP(n6800), .ZN(n6805));
   INVX0 U7372 (.INP(n6909), .ZN(n6908));
   INVX0 U7373 (.INP(n6881), .ZN(n6880));
   INVX0 U7374 (.INP(n7208), .ZN(n6909));
   INVX0 U7375 (.INP(n7006), .ZN(n6881));
   INVX0 U7376 (.INP(n6908), .ZN(n6906));
   INVX0 U7377 (.INP(n6908), .ZN(n6907));
   INVX0 U7378 (.INP(n6880), .ZN(n6879));
   INVX0 U7379 (.INP(n6880), .ZN(n6878));
   INVX0 U7380 (.INP(n6859), .ZN(n6852));
   INVX0 U7381 (.INP(n6859), .ZN(n6853));
   INVX0 U7382 (.INP(n6859), .ZN(n6858));
   INVX0 U7383 (.INP(n6859), .ZN(n6857));
   INVX0 U7384 (.INP(n6859), .ZN(n6854));
   INVX0 U7385 (.INP(n6859), .ZN(n6855));
   INVX0 U7386 (.INP(n6859), .ZN(n6856));
   INVX0 U7387 (.INP(n6988), .ZN(n6859));
   INVX0 U7388 (.INP(n6857), .ZN(n6842));
   INVX0 U7389 (.INP(n6852), .ZN(n6850));
   INVX0 U7390 (.INP(n6852), .ZN(n6851));
   INVX0 U7391 (.INP(n6853), .ZN(n6849));
   INVX0 U7392 (.INP(n6854), .ZN(n6847));
   INVX0 U7393 (.INP(n6854), .ZN(n6848));
   INVX0 U7394 (.INP(n6855), .ZN(n6845));
   INVX0 U7395 (.INP(n6855), .ZN(n6846));
   INVX0 U7396 (.INP(n6856), .ZN(n6843));
   INVX0 U7397 (.INP(n6856), .ZN(n6844));
   INVX0 U7398 (.INP(n6877), .ZN(n6869));
   INVX0 U7399 (.INP(n6877), .ZN(n6870));
   INVX0 U7400 (.INP(n6876), .ZN(n6875));
   INVX0 U7401 (.INP(n6876), .ZN(n6874));
   INVX0 U7402 (.INP(n6876), .ZN(n6871));
   INVX0 U7403 (.INP(n6876), .ZN(n6872));
   INVX0 U7404 (.INP(n6876), .ZN(n6873));
   INVX0 U7405 (.INP(n6989), .ZN(n6877));
   INVX0 U7406 (.INP(n6989), .ZN(n6876));
   INVX0 U7407 (.INP(n6874), .ZN(n6860));
   INVX0 U7408 (.INP(n6872), .ZN(n6863));
   INVX0 U7409 (.INP(n6873), .ZN(n6861));
   INVX0 U7410 (.INP(n6873), .ZN(n6862));
   INVX0 U7411 (.INP(n6869), .ZN(n6867));
   INVX0 U7412 (.INP(n6869), .ZN(n6868));
   INVX0 U7413 (.INP(n6870), .ZN(n6866));
   INVX0 U7414 (.INP(n6871), .ZN(n6864));
   INVX0 U7415 (.INP(n6871), .ZN(n6865));
   INVX0 U7416 (.INP(n6817), .ZN(n6808));
   INVX0 U7417 (.INP(n6815), .ZN(n6809));
   INVX0 U7418 (.INP(n6816), .ZN(n6810));
   INVX0 U7419 (.INP(n6816), .ZN(n6811));
   INVX0 U7420 (.INP(n6815), .ZN(n6812));
   INVX0 U7421 (.INP(n6815), .ZN(n6813));
   INVX0 U7422 (.INP(n2278), .ZN(n6814));
   INVX0 U7423 (.INP(n2278), .ZN(n6815));
   INVX0 U7424 (.INP(n2278), .ZN(n6816));
   INVX0 U7425 (.INP(n2278), .ZN(n6817));
   INVX0 U7426 (.INP(n6808), .ZN(n6818));
   INVX0 U7427 (.INP(n6808), .ZN(n6819));
   INVX0 U7428 (.INP(n6808), .ZN(n6820));
   INVX0 U7429 (.INP(n6808), .ZN(n6821));
   INVX0 U7430 (.INP(n6808), .ZN(n6822));
   INVX0 U7431 (.INP(n6808), .ZN(n6823));
   INVX0 U7432 (.INP(n6927), .ZN(n6824));
   INVX0 U7433 (.INP(n6927), .ZN(n6825));
   INVX0 U7434 (.INP(n6817), .ZN(n6927));
   INVX0 U7435 (.INP(n6815), .ZN(n6926));
   INVX0 U7436 (.INP(new_sboxw[25]), .ZN(n7592));
   NBUFFX2 U7437 (.INP(n7097), .Z(n7118));
   NBUFFX2 U7438 (.INP(n7097), .Z(n7116));
   NBUFFX2 U7439 (.INP(n7097), .Z(n7117));
   NBUFFX2 U7440 (.INP(n2295), .Z(n7093));
   NBUFFX2 U7441 (.INP(n2295), .Z(n7091));
   NBUFFX2 U7442 (.INP(n2295), .Z(n7092));
   NBUFFX2 U7443 (.INP(n2295), .Z(n7095));
   NBUFFX2 U7444 (.INP(n2295), .Z(n7096));
   NBUFFX2 U7445 (.INP(n2295), .Z(n7094));
   NBUFFX2 U7446 (.INP(n2295), .Z(n7097));
   INVX0 U7447 (.INP(new_sboxw[30]), .ZN(n7597));
   INVX0 U7448 (.INP(new_sboxw[10]), .ZN(n7606));
   INVX0 U7449 (.INP(new_sboxw[27]), .ZN(n7594));
   AND2X1 U7450 (.IN1(n7580), .IN2(n2214), .Q(n2295));
   INVX0 U7451 (.INP(new_sboxw[15]), .ZN(n7611));
   INVX0 U7452 (.INP(new_sboxw[12]), .ZN(n7608));
   INVX0 U7453 (.INP(new_sboxw[11]), .ZN(n7607));
   INVX0 U7454 (.INP(keylen), .ZN(n7622));
   INVX0 U7455 (.INP(n2957), .ZN(n7586));
   INVX0 U7456 (.INP(new_sboxw[18]), .ZN(n7601));
   INVX0 U7457 (.INP(new_sboxw[26]), .ZN(n7593));
   INVX0 U7458 (.INP(new_sboxw[31]), .ZN(n7598));
   INVX0 U7459 (.INP(new_sboxw[8]), .ZN(n7612));
   INVX0 U7460 (.INP(new_sboxw[20]), .ZN(n7603));
   INVX0 U7461 (.INP(new_sboxw[9]), .ZN(n7613));
   INVX0 U7462 (.INP(new_sboxw[19]), .ZN(n7602));
   INVX0 U7463 (.INP(new_sboxw[28]), .ZN(n7595));
   INVX0 U7464 (.INP(n7286), .ZN(n7285));
   INVX0 U7465 (.INP(n7288), .ZN(n7284));
   INVX0 U7466 (.INP(n6967), .ZN(n7229));
   INVX0 U7467 (.INP(n7230), .ZN(n7228));
   INVX0 U7468 (.INP(n6968), .ZN(n7205));
   INVX0 U7469 (.INP(n7206), .ZN(n7204));
   INVX0 U7470 (.INP(new_sboxw[21]), .ZN(n7604));
   INVX0 U7471 (.INP(n6925), .ZN(n7286));
   INVX0 U7472 (.INP(n2944), .ZN(n6943));
   INVX0 U7473 (.INP(n6943), .ZN(n6950));
   INVX0 U7474 (.INP(n6943), .ZN(n6951));
   INVX0 U7475 (.INP(n6943), .ZN(n6952));
   INVX0 U7476 (.INP(n6943), .ZN(n6953));
   INVX0 U7477 (.INP(n6943), .ZN(n6954));
   INVX0 U7478 (.INP(n6943), .ZN(n6955));
   INVX0 U7479 (.INP(n3395), .ZN(n6956));
   INVX0 U7480 (.INP(n6956), .ZN(n6961));
   INVX0 U7481 (.INP(n6956), .ZN(n6962));
   INVX0 U7482 (.INP(n6956), .ZN(n6963));
   INVX0 U7483 (.INP(n6956), .ZN(n6964));
   INVX0 U7484 (.INP(n6956), .ZN(n6965));
   NOR2X0 U7485 (.IN1(n7580), .IN2(n6964), .QN(n3396));
   INVX0 U7486 (.INP(new_sboxw[4]), .ZN(n7618));
   INVX0 U7487 (.INP(new_sboxw[3]), .ZN(n7617));
   INVX0 U7488 (.INP(new_sboxw[2]), .ZN(n7616));
   INVX0 U7489 (.INP(new_sboxw[1]), .ZN(n7615));
   INVX0 U7490 (.INP(new_sboxw[7]), .ZN(n7621));
   INVX0 U7491 (.INP(new_sboxw[6]), .ZN(n7620));
   INVX0 U7492 (.INP(new_sboxw[5]), .ZN(n7619));
   NOR2X0 U7493 (.IN1(n7622), .IN2(n6814), .QN(n2297));
   INVX0 U7494 (.INP(new_sboxw[14]), .ZN(n7610));
   INVX0 U7495 (.INP(new_sboxw[0]), .ZN(n7614));
   INVX0 U7496 (.INP(new_sboxw[13]), .ZN(n7609));
   INVX0 U7497 (.INP(new_sboxw[24]), .ZN(n7591));
   INVX0 U7498 (.INP(n2948), .ZN(n7589));
   INVX0 U7499 (.INP(new_sboxw[17]), .ZN(n7600));
   INVX0 U7500 (.INP(n7010), .ZN(n7011));
   INVX0 U7501 (.INP(n7005), .ZN(n7006));
   INVX0 U7502 (.INP(n7021), .ZN(n7022));
   INVX0 U7503 (.INP(n6966), .ZN(n7312));
   INVX0 U7504 (.INP(n6966), .ZN(n7311));
   INVX0 U7505 (.INP(n7310), .ZN(n7309));
   INVX0 U7506 (.INP(n6966), .ZN(n7305));
   INVX0 U7507 (.INP(n6966), .ZN(n7306));
   INVX0 U7508 (.INP(n7310), .ZN(n7307));
   INVX0 U7509 (.INP(n7310), .ZN(n7308));
   INVX0 U7510 (.INP(n7310), .ZN(n7300));
   INVX0 U7511 (.INP(n6966), .ZN(n7301));
   INVX0 U7512 (.INP(n7310), .ZN(n7302));
   INVX0 U7513 (.INP(n6966), .ZN(n7303));
   INVX0 U7514 (.INP(n7310), .ZN(n7304));
   INVX0 U7515 (.INP(n6966), .ZN(n7295));
   INVX0 U7516 (.INP(n7310), .ZN(n7296));
   INVX0 U7517 (.INP(n7310), .ZN(n7297));
   INVX0 U7518 (.INP(n7310), .ZN(n7298));
   INVX0 U7519 (.INP(n7310), .ZN(n7299));
   INVX0 U7520 (.INP(n7310), .ZN(n7290));
   INVX0 U7521 (.INP(n7310), .ZN(n7291));
   INVX0 U7522 (.INP(n7310), .ZN(n7292));
   INVX0 U7523 (.INP(n6966), .ZN(n7293));
   INVX0 U7524 (.INP(n7310), .ZN(n7294));
   AOI21X1 U7525 (.IN1(n3401), .IN2(n7581), .IN3(n3405), .QN(n2944));
   INVX0 U7526 (.INP(n7234), .ZN(n6967));
   INVX0 U7527 (.INP(n6993), .ZN(n7234));
   INVX0 U7528 (.INP(n7210), .ZN(n6968));
   INVX0 U7529 (.INP(n6991), .ZN(n7210));
   INVX0 U7530 (.INP(n2283), .ZN(n6969));
   INVX0 U7531 (.INP(n2283), .ZN(n6970));
   INVX0 U7532 (.INP(n2283), .ZN(n7266));
   INVX0 U7533 (.INP(n7015), .ZN(n7017));
   INVX0 U7534 (.INP(n7015), .ZN(n7016));
   INVX0 U7535 (.INP(n7265), .ZN(n7015));
   INVX0 U7536 (.INP(n7264), .ZN(n7251));
   INVX0 U7537 (.INP(n7260), .ZN(n7259));
   INVX0 U7538 (.INP(n7260), .ZN(n7258));
   INVX0 U7539 (.INP(n7261), .ZN(n7256));
   INVX0 U7540 (.INP(n7261), .ZN(n7257));
   INVX0 U7541 (.INP(n7262), .ZN(n7254));
   INVX0 U7542 (.INP(n7262), .ZN(n7255));
   INVX0 U7543 (.INP(n7263), .ZN(n7252));
   INVX0 U7544 (.INP(n7263), .ZN(n7253));
   INVX0 U7545 (.INP(n7287), .ZN(n7021));
   INVX0 U7546 (.INP(n7231), .ZN(n7010));
   INVX0 U7547 (.INP(n7207), .ZN(n7005));
   INVX0 U7548 (.INP(n7165), .ZN(n6971));
   INVX0 U7549 (.INP(n7165), .ZN(n6972));
   INVX0 U7550 (.INP(n7152), .ZN(n7158));
   INVX0 U7551 (.INP(n7153), .ZN(n7159));
   INVX0 U7552 (.INP(n6994), .ZN(n6996));
   INVX0 U7553 (.INP(n6994), .ZN(n6995));
   INVX0 U7554 (.INP(n7163), .ZN(n6994));
   INVX0 U7555 (.INP(n7160), .ZN(n7152));
   INVX0 U7556 (.INP(n7160), .ZN(n7153));
   INVX0 U7557 (.INP(n7161), .ZN(n7150));
   INVX0 U7558 (.INP(n7161), .ZN(n7151));
   INVX0 U7559 (.INP(n7162), .ZN(n7148));
   INVX0 U7560 (.INP(n7162), .ZN(n7149));
   INVX0 U7561 (.INP(n7158), .ZN(n7156));
   INVX0 U7562 (.INP(n7158), .ZN(n7157));
   INVX0 U7563 (.INP(n7159), .ZN(n7154));
   INVX0 U7564 (.INP(n7159), .ZN(n7155));
   INVX0 U7565 (.INP(n6995), .ZN(n7147));
   INVX0 U7566 (.INP(n7281), .ZN(n6973));
   INVX0 U7567 (.INP(n7281), .ZN(n6974));
   INVX0 U7568 (.INP(n7282), .ZN(n7274));
   INVX0 U7569 (.INP(n7282), .ZN(n7275));
   INVX0 U7570 (.INP(n7281), .ZN(n7280));
   INVX0 U7571 (.INP(n7281), .ZN(n7278));
   INVX0 U7572 (.INP(n7018), .ZN(n7020));
   INVX0 U7573 (.INP(n7018), .ZN(n7019));
   INVX0 U7574 (.INP(n7279), .ZN(n7018));
   INVX0 U7575 (.INP(n7277), .ZN(n7268));
   INVX0 U7576 (.INP(n7276), .ZN(n7269));
   INVX0 U7577 (.INP(n7276), .ZN(n7270));
   INVX0 U7578 (.INP(n7274), .ZN(n7273));
   INVX0 U7579 (.INP(n7275), .ZN(n7271));
   INVX0 U7580 (.INP(n7275), .ZN(n7272));
   INVX0 U7581 (.INP(n7278), .ZN(n7267));
   INVX0 U7582 (.INP(n7225), .ZN(n6975));
   INVX0 U7583 (.INP(n7225), .ZN(n6976));
   INVX0 U7584 (.INP(n7226), .ZN(n7218));
   INVX0 U7585 (.INP(n7226), .ZN(n7219));
   INVX0 U7586 (.INP(n7225), .ZN(n7224));
   INVX0 U7587 (.INP(n7225), .ZN(n7222));
   INVX0 U7588 (.INP(n7007), .ZN(n7009));
   INVX0 U7589 (.INP(n7007), .ZN(n7008));
   INVX0 U7590 (.INP(n7223), .ZN(n7007));
   INVX0 U7591 (.INP(n7221), .ZN(n7212));
   INVX0 U7592 (.INP(n7221), .ZN(n7213));
   INVX0 U7593 (.INP(n7220), .ZN(n7214));
   INVX0 U7594 (.INP(n7218), .ZN(n7217));
   INVX0 U7595 (.INP(n7219), .ZN(n7215));
   INVX0 U7596 (.INP(n7219), .ZN(n7216));
   INVX0 U7597 (.INP(n7222), .ZN(n7211));
   INVX0 U7598 (.INP(n7201), .ZN(n6977));
   INVX0 U7599 (.INP(n7201), .ZN(n6978));
   INVX0 U7600 (.INP(n7202), .ZN(n7194));
   INVX0 U7601 (.INP(n7202), .ZN(n7195));
   INVX0 U7602 (.INP(n7201), .ZN(n7200));
   INVX0 U7603 (.INP(n7201), .ZN(n7198));
   INVX0 U7604 (.INP(n7002), .ZN(n7004));
   INVX0 U7605 (.INP(n7002), .ZN(n7003));
   INVX0 U7606 (.INP(n7199), .ZN(n7002));
   INVX0 U7607 (.INP(n7197), .ZN(n7188));
   INVX0 U7608 (.INP(n7197), .ZN(n7189));
   INVX0 U7609 (.INP(n7196), .ZN(n7190));
   INVX0 U7610 (.INP(n7194), .ZN(n7193));
   INVX0 U7611 (.INP(n7195), .ZN(n7191));
   INVX0 U7612 (.INP(n7195), .ZN(n7192));
   INVX0 U7613 (.INP(n7198), .ZN(n7187));
   INVX0 U7614 (.INP(n7180), .ZN(n6979));
   INVX0 U7615 (.INP(n7180), .ZN(n6980));
   INVX0 U7616 (.INP(n7181), .ZN(n7173));
   INVX0 U7617 (.INP(n7181), .ZN(n7174));
   INVX0 U7618 (.INP(n7180), .ZN(n7179));
   INVX0 U7619 (.INP(n7180), .ZN(n7177));
   INVX0 U7620 (.INP(n6997), .ZN(n6999));
   INVX0 U7621 (.INP(n6997), .ZN(n6998));
   INVX0 U7622 (.INP(n7178), .ZN(n6997));
   INVX0 U7623 (.INP(n7176), .ZN(n7167));
   INVX0 U7624 (.INP(n7176), .ZN(n7168));
   INVX0 U7625 (.INP(n7175), .ZN(n7169));
   INVX0 U7626 (.INP(n7173), .ZN(n7172));
   INVX0 U7627 (.INP(n7174), .ZN(n7170));
   INVX0 U7628 (.INP(n7174), .ZN(n7171));
   INVX0 U7629 (.INP(n7177), .ZN(n7166));
   INVX0 U7630 (.INP(new_sboxw[16]), .ZN(n7599));
   INVX0 U7631 (.INP(new_sboxw[29]), .ZN(n7596));
   INVX0 U7632 (.INP(n7311), .ZN(n7310));
   INVX0 U7633 (.INP(n7186), .ZN(n6981));
   INVX0 U7634 (.INP(n7186), .ZN(n6982));
   INVX0 U7635 (.INP(n6986), .ZN(n6983));
   INVX0 U7636 (.INP(n7001), .ZN(n6984));
   INVX0 U7637 (.INP(n7001), .ZN(n6985));
   INVX0 U7638 (.INP(n6981), .ZN(n6986));
   INVX0 U7639 (.INP(n6982), .ZN(n6987));
   INVX0 U7640 (.INP(n7183), .ZN(n7000));
   INVX0 U7641 (.INP(n7184), .ZN(n7183));
   INVX0 U7642 (.INP(n7000), .ZN(n7001));
   INVX0 U7643 (.INP(n2283), .ZN(n7265));
   INVX0 U7644 (.INP(n2283), .ZN(n7264));
   INVX0 U7645 (.INP(n2283), .ZN(n7263));
   INVX0 U7646 (.INP(n2283), .ZN(n7262));
   INVX0 U7647 (.INP(n2283), .ZN(n7261));
   INVX0 U7648 (.INP(n2283), .ZN(n7260));
   NAND2X0 U7649 (.IN1(n2935), .IN2(n2931), .QN(n2283));
   NAND2X1 U7650 (.IN1(n2935), .IN2(n2933), .QN(n2284));
   INVX0 U7651 (.INP(n7249), .ZN(n7012));
   INVX0 U7652 (.INP(n7244), .ZN(n7243));
   INVX0 U7653 (.INP(n7248), .ZN(n7235));
   INVX0 U7654 (.INP(n7248), .ZN(n7236));
   INVX0 U7655 (.INP(n7247), .ZN(n7237));
   INVX0 U7656 (.INP(n7247), .ZN(n7238));
   INVX0 U7657 (.INP(n7246), .ZN(n7239));
   INVX0 U7658 (.INP(n7246), .ZN(n7240));
   INVX0 U7659 (.INP(n7245), .ZN(n7241));
   INVX0 U7660 (.INP(n7245), .ZN(n7242));
   INVX0 U7661 (.INP(n2284), .ZN(n7249));
   INVX0 U7662 (.INP(n2284), .ZN(n7250));
   INVX0 U7663 (.INP(n2284), .ZN(n7248));
   INVX0 U7664 (.INP(n2284), .ZN(n7247));
   INVX0 U7665 (.INP(n2284), .ZN(n7246));
   INVX0 U7666 (.INP(n2284), .ZN(n7245));
   INVX0 U7667 (.INP(n2284), .ZN(n7244));
   INVX0 U7668 (.INP(n7012), .ZN(n7014));
   INVX0 U7669 (.INP(n7012), .ZN(n7013));
   NOR2X0 U7670 (.IN1(round_ctr_reg[2]), .IN2(n2213), .QN(n3417));
   INVX0 U7671 (.INP(n7289), .ZN(n7288));
   INVX0 U7672 (.INP(n7289), .ZN(n7287));
   INVX0 U7673 (.INP(n6990), .ZN(n7289));
   INVX0 U7674 (.INP(n7233), .ZN(n7231));
   INVX0 U7675 (.INP(n7233), .ZN(n7230));
   INVX0 U7676 (.INP(n7233), .ZN(n7232));
   INVX0 U7677 (.INP(n6993), .ZN(n7233));
   INVX0 U7678 (.INP(n7209), .ZN(n7208));
   INVX0 U7679 (.INP(n7209), .ZN(n7207));
   INVX0 U7680 (.INP(n7209), .ZN(n7206));
   INVX0 U7681 (.INP(n6991), .ZN(n7209));
   INVX0 U7682 (.INP(n7165), .ZN(n7164));
   INVX0 U7683 (.INP(n7165), .ZN(n7163));
   INVX0 U7684 (.INP(n7165), .ZN(n7162));
   INVX0 U7685 (.INP(n7165), .ZN(n7161));
   INVX0 U7686 (.INP(n7165), .ZN(n7160));
   INVX0 U7687 (.INP(n6992), .ZN(n7165));
   INVX0 U7688 (.INP(n7283), .ZN(n7281));
   INVX0 U7689 (.INP(n7281), .ZN(n7279));
   INVX0 U7690 (.INP(n7283), .ZN(n7282));
   INVX0 U7691 (.INP(n7281), .ZN(n7276));
   INVX0 U7692 (.INP(n7281), .ZN(n7277));
   INVX0 U7693 (.INP(n7227), .ZN(n7225));
   INVX0 U7694 (.INP(n7225), .ZN(n7223));
   INVX0 U7695 (.INP(n7227), .ZN(n7226));
   INVX0 U7696 (.INP(n7225), .ZN(n7220));
   INVX0 U7697 (.INP(n7225), .ZN(n7221));
   INVX0 U7698 (.INP(n7203), .ZN(n7201));
   INVX0 U7699 (.INP(n7201), .ZN(n7199));
   INVX0 U7700 (.INP(n7203), .ZN(n7202));
   INVX0 U7701 (.INP(n7201), .ZN(n7196));
   INVX0 U7702 (.INP(n7201), .ZN(n7197));
   INVX0 U7703 (.INP(n7182), .ZN(n7180));
   INVX0 U7704 (.INP(n7180), .ZN(n7178));
   INVX0 U7705 (.INP(n7182), .ZN(n7181));
   INVX0 U7706 (.INP(n7180), .ZN(n7175));
   INVX0 U7707 (.INP(n7180), .ZN(n7176));
   INVX0 U7708 (.INP(n3397), .ZN(n7580));
   NOR2X0 U7709 (.IN1(n3410), .IN2(n2941), .QN(n3411));
   INVX0 U7710 (.INP(n2282), .ZN(n7283));
   INVX0 U7711 (.INP(n2286), .ZN(n7227));
   INVX0 U7712 (.INP(n2288), .ZN(n7203));
   NOR2X0 U7713 (.IN1(n2212), .IN2(round_ctr_reg[2]), .QN(n2936));
   NOR2X0 U7714 (.IN1(n2941), .IN2(round_ctr_reg[0]), .QN(n2931));
   NAND2X0 U7715 (.IN1(n2243), .IN2(key_mem_ctrl_reg[1]), .QN(n2941));
   INVX0 U7716 (.INP(n2289), .ZN(n7186));
   INVX0 U7717 (.INP(n7186), .ZN(n7184));
   INVX0 U7718 (.INP(n7186), .ZN(n7185));
   INVX0 U7719 (.INP(n2290), .ZN(n7182));
   NOR2X0 U7720 (.IN1(n2214), .IN2(n2941), .QN(n2933));
   NAND2X0 U7721 (.IN1(n3407), .IN2(n2214), .QN(n3403));
   NOR2X0 U7722 (.IN1(n6966), .IN2(n7622), .QN(n3395));
   NOR2X0 U7723 (.IN1(n3406), .IN2(n2941), .QN(n2278));
   NOR2X0 U7724 (.IN1(n6966), .IN2(n6944), .QN(n2945));
   NAND2X0 U7725 (.IN1(round_ctr_reg[0]), .IN2(n3407), .QN(n3406));
   NAND3X0 U7726 (.IN1(n2243), .IN2(n2242), .IN3(init), .QN(n3408));
   assign clk_buf_net0 = clk;
   assign clk_buf_net1 = clk_buf_net0;
   assign clk_buf_net2 = clk_buf_net1;
   assign clk_buf_net3 = clk_buf_net2;
   assign clk_buf_net4 = clk_buf_net3;
   assign clk_buf_net5 = clk_buf_net4;
   assign clk_buf_net6 = clk_buf_net5;
   assign clk_buf_net7 = clk_buf_net6;
   assign test_se_buf_net0 = test_se;
   assign test_se_buf_net1 = test_se_buf_net0;
   assign test_se_buf_net2 = test_se_buf_net1;
   assign test_se_buf_net3 = test_se_buf_net2;
   assign test_se_buf_net4 = test_se_buf_net3;
   assign test_se_buf_net5 = test_se_buf_net4;
   assign test_se_buf_net6 = test_se_buf_net5;
   assign test_se_buf_net7 = test_se_buf_net6;
endmodule

module aes_sbox (sboxw, new_sboxw);
input [31:0] sboxw;
output [31:0] new_sboxw;
wire n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
       n200, n201, n202, n203, n204, n206, n207, n208, n209, n210, n211, n212, n213, n214
       , n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
       n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241
       , n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
       n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268
       , n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
       n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295
       , n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
       n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322
       , n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
       n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350
       , n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
       n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377
       , n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
       n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404
       , n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
       n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431
       , n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
       n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458
       , n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
       n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485
       , n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
       n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512
       , n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
       n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539
       , n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
       n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n565, n566, n567
       , n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
       n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594
       , n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
       n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621
       , n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
       n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648
       , n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, 
       n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675
       , n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
       n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702
       , n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
       n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729
       , n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
       n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756
       , n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, 
       n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783
       , n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, 
       n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810
       , n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
       n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837
       , n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, 
       n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864
       , n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, 
       n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891
       , n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, 
       n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918
       , n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
       n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945
       , n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, 
       n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972
       , n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, 
       n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999
       , n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
       n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022
       , n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
       n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045
       , n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, 
       n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068
       , n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
       n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091
       , n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
       n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114
       , n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, 
       n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137
       , n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
       n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160
       , n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, 
       n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183
       , n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
       n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206
       , n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, 
       n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229
       , n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, 
       n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252
       , n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
       n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275
       , n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, 
       n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298
       , n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
       n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321
       , n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
       n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344
       , n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
       n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367
       , n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
       n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390
       , n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, 
       n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413
       , n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
       n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436
       , n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
       n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459
       , n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, 
       n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482
       , n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, 
       n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505
       , n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, 
       n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528
       , n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1, 
       n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, 
       n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
       , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
       n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69
       , n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, 
       n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
       n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115
       , n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, 
       n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142
       , n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
       n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169
       , n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
       n183, n184, n185, n205, n323, n564, n1540, n1541, n1542, n1543, n1544, n1545, n1546
       , n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, 
       n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569
       , n1570, n1571;
   AO22X1 U753 (.IN1(sboxw[15]), .IN2(n186), .IN3(n187), .IN4(n134), .Q(new_sboxw[9]));
   AO222X1 U754 (.IN1(n188), .IN2(n189), .IN3(n190), .IN4(n191), .IN5(n192), .IN6(n135), .
          Q(n187));
   NAND4X0 U755 (.IN1(n193), .IN2(n194), .IN3(n195), .IN4(n196), .QN(n192));
   OA221X1 U756 (.IN1(n197), .IN2(n159), .IN3(n198), .IN4(n143), .IN5(n199), .Q(n196));
   AOI22X1 U757 (.IN1(n173), .IN2(n200), .IN3(n27), .IN4(n202), .QN(n199));
   OA22X1 U758 (.IN1(n203), .IN2(n43), .IN3(n204), .IN4(n137), .Q(n195));
   OA22X1 U759 (.IN1(n177), .IN2(n152), .IN3(n38), .IN4(n147), .Q(n203));
   NAND3X0 U760 (.IN1(n43), .IN2(n177), .IN3(n206), .QN(n193));
   NAND4X0 U761 (.IN1(n207), .IN2(n208), .IN3(n209), .IN4(n210), .QN(n191));
   OA222X1 U762 (.IN1(n175), .IN2(n152), .IN3(n211), .IN4(n146), .IN5(n162), .IN6(n173), .
          Q(n210));
   OA22X1 U763 (.IN1(n204), .IN2(n212), .IN3(n150), .IN4(n177), .Q(n209));
   NAND4X0 U764 (.IN1(n213), .IN2(n214), .IN3(n215), .IN4(n216), .QN(n189));
   OA222X1 U765 (.IN1(n211), .IN2(n163), .IN3(n150), .IN4(n175), .IN5(n152), .IN6(n3), .Q(
          n216));
   OA22X1 U766 (.IN1(n177), .IN2(n165), .IN3(n38), .IN4(n217), .Q(n215));
   AO221X1 U767 (.IN1(n188), .IN2(n218), .IN3(n219), .IN4(n135), .IN5(n220), .Q(n186));
   AO22X1 U768 (.IN1(n190), .IN2(n221), .IN3(n222), .IN4(n223), .Q(n220));
   NAND4X0 U769 (.IN1(n224), .IN2(n225), .IN3(n226), .IN4(n227), .QN(n221));
   OA22X1 U770 (.IN1(n37), .IN2(n152), .IN3(n148), .IN4(n3), .Q(n227));
   AO222X1 U771 (.IN1(n229), .IN2(n230), .IN3(n9), .IN4(n231), .IN5(n232), .IN6(n43), .Q(
          n219));
   NAND3X0 U772 (.IN1(n233), .IN2(n234), .IN3(n235), .QN(n232));
   OA222X1 U773 (.IN1(n172), .IN2(n236), .IN3(n173), .IN4(n237), .IN5(n41), .IN6(n145), .Q(
          n235));
   OA22X1 U774 (.IN1(n211), .IN2(n161), .IN3(n27), .IN4(n158), .Q(n233));
   NAND3X0 U775 (.IN1(n238), .IN2(n239), .IN3(n240), .QN(n231));
   AO221X1 U776 (.IN1(n241), .IN2(n177), .IN3(n242), .IN4(n173), .IN5(n243), .Q(n230));
   AO22X1 U777 (.IN1(n18), .IN2(n244), .IN3(n245), .IN4(n175), .Q(n243));
   OA222X1 U778 (.IN1(n146), .IN2(n173), .IN3(n248), .IN4(n177), .IN5(n212), .IN6(n174), .
          Q(n247));
   OA222X1 U779 (.IN1(n163), .IN2(n3), .IN3(n18), .IN4(n162), .IN5(n204), .IN6(n152), .Q(
          n246));
   AO22X1 U780 (.IN1(sboxw[15]), .IN2(n251), .IN3(n252), .IN4(n134), .Q(new_sboxw[8]));
   AO22X1 U781 (.IN1(n253), .IN2(n135), .IN3(sboxw[14]), .IN4(n254), .Q(n252));
   NAND4X0 U782 (.IN1(n255), .IN2(n144), .IN3(n256), .IN4(n257), .QN(n254));
   AOI222X1 U783 (.IN1(n9), .IN2(n258), .IN3(n259), .IN4(n43), .IN5(n260), .IN6(n42), .QN(
          n257));
   AO221X1 U784 (.IN1(n242), .IN2(n261), .IN3(n204), .IN4(n245), .IN5(n262), .Q(n259));
   NAND4X0 U785 (.IN1(n238), .IN2(n158), .IN3(n263), .IN4(n264), .QN(n258));
   OA222X1 U786 (.IN1(n159), .IN2(n177), .IN3(n173), .IN4(n265), .IN5(n146), .IN6(n3), .Q(
          n264));
   NAND3X0 U787 (.IN1(n37), .IN2(n20), .IN3(n271), .QN(n255));
   NAND4X0 U788 (.IN1(n272), .IN2(n273), .IN3(n274), .IN4(n275), .QN(n253));
   AOI222X1 U789 (.IN1(n9), .IN2(n276), .IN3(n277), .IN4(n175), .IN5(n260), .IN6(n176), .
          QN(n275));
   NAND4X0 U790 (.IN1(n278), .IN2(n239), .IN3(n279), .IN4(n280), .QN(n276));
   OA222X1 U791 (.IN1(n29), .IN2(n147), .IN3(n146), .IN4(n175), .IN5(n281), .IN6(n162), .Q(
          n280));
   NAND3X0 U792 (.IN1(n154), .IN2(n174), .IN3(n271), .QN(n272));
   AO222X1 U793 (.IN1(sboxw[14]), .IN2(n283), .IN3(n188), .IN4(n284), .IN5(n285), .IN6(
          n135), .Q(n251));
   AO221X1 U794 (.IN1(n286), .IN2(n287), .IN3(n288), .IN4(n43), .IN5(n289), .Q(n285));
   AO222X1 U795 (.IN1(n290), .IN2(n176), .IN3(n291), .IN4(n19), .IN5(n281), .IN6(n223), .Q(
          n289));
   OAI221X1 U796 (.IN1(n162), .IN2(n204), .IN3(n158), .IN4(n27), .IN5(n225), .QN(n288));
   AO221X1 U797 (.IN1(n241), .IN2(n174), .IN3(n245), .IN4(n177), .IN5(n293), .Q(n287));
   AO221X1 U798 (.IN1(n281), .IN2(n206), .IN3(n242), .IN4(n261), .IN5(n149), .Q(n284));
   AO22X1 U799 (.IN1(n18), .IN2(n172), .IN3(n19), .IN4(n3), .Q(n261));
   AO221X1 U800 (.IN1(n294), .IN2(n286), .IN3(n9), .IN4(n295), .IN5(n269), .Q(n283));
   NAND3X0 U801 (.IN1(n296), .IN2(n297), .IN3(n298), .QN(n295));
   AOI221X1 U802 (.IN1(n204), .IN2(n299), .IN3(n175), .IN4(n300), .IN5(n301), .QN(n298));
   OA22X1 U803 (.IN1(n281), .IN2(n217), .IN3(n177), .IN4(n162), .Q(n296));
   AO222X1 U804 (.IN1(n302), .IN2(n303), .IN3(n304), .IN4(n305), .IN5(n306), .IN6(n178), .
          Q(new_sboxw[7]));
   AO222X1 U805 (.IN1(n307), .IN2(n308), .IN3(n309), .IN4(n310), .IN5(n311), .IN6(n179), .
          Q(n306));
   NAND4X0 U806 (.IN1(n312), .IN2(n313), .IN3(n314), .IN4(n315), .QN(n311));
   AOI222X1 U807 (.IN1(n316), .IN2(n12), .IN3(n317), .IN4(n1569), .IN5(n8), .IN6(n318), .
          QN(n315));
   NAND4X0 U808 (.IN1(n319), .IN2(n1543), .IN3(n320), .IN4(n321), .QN(n318));
   OA22X1 U809 (.IN1(n35), .IN2(n324), .IN3(n1552), .IN4(n325), .Q(n314));
   NAND3X0 U810 (.IN1(n1567), .IN2(n1564), .IN3(n327), .QN(n312));
   NAND4X0 U811 (.IN1(n1565), .IN2(n328), .IN3(n329), .IN4(n330), .QN(n310));
   OA222X1 U812 (.IN1(n331), .IN2(n1551), .IN3(n1571), .IN4(n332), .IN5(n36), .IN6(n1549)
          , .Q(n330));
   AND2X1 U813 (.IN1(n1556), .IN2(n333), .Q(n329));
   NAND4X0 U814 (.IN1(n335), .IN2(n336), .IN3(n337), .IN4(n338), .QN(n308));
   OA22X1 U815 (.IN1(n339), .IN2(n1571), .IN3(n1570), .IN4(n1556), .Q(n338));
   NAND3X0 U816 (.IN1(n35), .IN2(n16), .IN3(n340), .QN(n337));
   NAND3X0 U817 (.IN1(n17), .IN2(n341), .IN3(n342), .QN(n335));
   NAND4X0 U818 (.IN1(n343), .IN2(n180), .IN3(n344), .IN4(n345), .QN(n305));
   OA222X1 U819 (.IN1(n183), .IN2(n346), .IN3(n347), .IN4(n40), .IN5(n7), .IN6(n184), .Q(
          n345));
   AND3X1 U820 (.IN1(n348), .IN2(n1550), .IN3(n328), .Q(n347));
   OA22X1 U821 (.IN1(n350), .IN2(n323), .IN3(n8), .IN4(n351), .Q(n344));
   AND3X1 U822 (.IN1(n352), .IN2(n353), .IN3(n354), .Q(n351));
   NOR3X0 U823 (.IN1(n355), .IN2(n356), .IN3(n357), .QN(n350));
   OA221X1 U824 (.IN1(n1551), .IN2(n325), .IN3(n17), .IN4(n362), .IN5(n363), .Q(n361));
   OA22X1 U825 (.IN1(n331), .IN2(n1540), .IN3(n323), .IN4(n1569), .Q(n362));
   NAND3X0 U827 (.IN1(n367), .IN2(n368), .IN3(n369), .QN(n364));
   OA222X1 U828 (.IN1(n370), .IN2(n1560), .IN3(n36), .IN4(n332), .IN5(n1570), .IN6(n1549)
          , .Q(n369));
   AO222X1 U830 (.IN1(n373), .IN2(n374), .IN3(n375), .IN4(n376), .IN5(sboxw[6]), .IN6(n377)
          , .Q(n372));
   AO221X1 U831 (.IN1(n8), .IN2(n378), .IN3(n379), .IN4(n40), .IN5(n380), .Q(n377));
   AO22X1 U832 (.IN1(n331), .IN2(n381), .IN3(n317), .IN4(n36), .Q(n380));
   OA221X1 U833 (.IN1(n342), .IN2(n1546), .IN3(n15), .IN4(n384), .IN5(n385), .Q(n383));
   NAND3X0 U834 (.IN1(n1566), .IN2(n1553), .IN3(n370), .QN(n385));
   OA222X1 U835 (.IN1(n388), .IN2(n1552), .IN3(n1555), .IN4(n1), .IN5(n1561), .IN6(n1569)
          , .Q(n382));
   NAND3X0 U836 (.IN1(n389), .IN2(n353), .IN3(n390), .QN(n378));
   NAND4X0 U837 (.IN1(n392), .IN2(n393), .IN3(n394), .IN4(n395), .QN(n376));
   OA222X1 U838 (.IN1(n12), .IN2(n1549), .IN3(n396), .IN4(n397), .IN5(n39), .IN6(n1546), .
          Q(n395));
   OR2X1 U839 (.IN1(n398), .IN2(n15), .Q(n394));
   NAND4X0 U840 (.IN1(n333), .IN2(n1549), .IN3(n399), .IN4(n400), .QN(n374));
   OA222X1 U841 (.IN1(sboxw[1]), .IN2(n1552), .IN3(n1567), .IN4(n1545), .IN5(n342), .IN6(
          n1555), .Q(n400));
   OA22X1 U842 (.IN1(n391), .IN2(n401), .IN3(n1569), .IN4(n1556), .Q(n399));
   AO221X1 U843 (.IN1(n307), .IN2(n402), .IN3(n403), .IN4(n179), .IN5(n404), .Q(n371));
   AO22X1 U844 (.IN1(n405), .IN2(sboxw[6]), .IN3(n309), .IN4(n406), .Q(n404));
   OA221X1 U845 (.IN1(n15), .IN2(n1546), .IN3(n1), .IN4(n1542), .IN5(n409), .Q(n408));
   AOI222X1 U846 (.IN1(n1553), .IN2(n410), .IN3(n39), .IN4(n322), .IN5(n411), .IN6(n396), .
          QN(n407));
   OA221X1 U847 (.IN1(n414), .IN2(n183), .IN3(n415), .IN4(n1540), .IN5(n1559), .Q(n413));
   AND2X1 U848 (.IN1(n1543), .IN2(n416), .Q(n414));
   OA222X1 U849 (.IN1(n417), .IN2(n1557), .IN3(n418), .IN4(n40), .IN5(n8), .IN6(n419), .Q(
          n412));
   OA22X1 U850 (.IN1(n417), .IN2(n1552), .IN3(sboxw[3]), .IN4(n370), .Q(n419));
   NAND4X0 U851 (.IN1(n420), .IN2(n421), .IN3(n422), .IN4(n423), .QN(n402));
   OR2X1 U852 (.IN1(n1561), .IN2(n388), .Q(n421));
   AO222X1 U854 (.IN1(n366), .IN2(n427), .IN3(n428), .IN4(n40), .IN5(n8), .IN6(n429), .Q(
          n426));
   NAND4X0 U855 (.IN1(n346), .IN2(n321), .IN3(n328), .IN4(n430), .QN(n429));
   OA221X1 U856 (.IN1(n1), .IN2(n1560), .IN3(n431), .IN4(n1568), .IN5(n1562), .Q(n430));
   NAND3X0 U857 (.IN1(n1544), .IN2(n320), .IN3(n434), .QN(n428));
   AO221X1 U858 (.IN1(n17), .IN2(n1568), .IN3(n1571), .IN4(n1553), .IN5(n1564), .Q(n427)
          );
   AO22X1 U859 (.IN1(n435), .IN2(n179), .IN3(sboxw[6]), .IN4(n436), .Q(n425));
   AO221X1 U860 (.IN1(n366), .IN2(n437), .IN3(n8), .IN4(n438), .IN5(n439), .Q(n436));
   AO22X1 U861 (.IN1(n440), .IN2(n15), .IN3(n441), .IN4(n327), .Q(n439));
   NAND4X0 U862 (.IN1(n353), .IN2(n442), .IN3(n443), .IN4(n444), .QN(n438));
   OA221X1 U863 (.IN1(n39), .IN2(n1556), .IN3(n396), .IN4(n1549), .IN5(n445), .Q(n444));
   AO222X1 U864 (.IN1(n396), .IN2(n391), .IN3(n35), .IN4(n447), .IN5(n411), .IN6(n1570), .
          Q(n437));
   NAND4X0 U865 (.IN1(n1554), .IN2(n442), .IN3(n448), .IN4(n449), .QN(n435));
   OA221X1 U866 (.IN1(n450), .IN2(n40), .IN3(n8), .IN4(n451), .IN5(n452), .Q(n449));
   OA22X1 U867 (.IN1(n453), .IN2(n183), .IN3(n396), .IN4(n1556), .Q(n452));
   AND3X1 U868 (.IN1(n1544), .IN2(n1561), .IN3(n416), .Q(n453));
   NAND4X0 U869 (.IN1(n313), .IN2(n336), .IN3(n456), .IN4(n457), .QN(n424));
   OA222X1 U870 (.IN1(n458), .IN2(n40), .IN3(n8), .IN4(n459), .IN5(n184), .IN6(n1), .Q(
          n457));
   OA22X1 U871 (.IN1(n1545), .IN2(sboxw[1]), .IN3(n1558), .IN4(n342), .Q(n367));
   OA221X1 U872 (.IN1(n39), .IN2(n1561), .IN3(n36), .IN4(n1551), .IN5(n461), .Q(n458));
   OA22X1 U873 (.IN1(n183), .IN2(n462), .IN3(n463), .IN4(n323), .Q(n456));
   NAND3X0 U874 (.IN1(n464), .IN2(n1), .IN3(n391), .QN(n313));
   AO22X1 U875 (.IN1(n465), .IN2(n178), .IN3(sboxw[7]), .IN4(n466), .Q(new_sboxw[4]));
   AO222X1 U876 (.IN1(n373), .IN2(n467), .IN3(n375), .IN4(n468), .IN5(sboxw[6]), .IN6(n469)
          , .Q(n466));
   OAI222X1 U877 (.IN1(n470), .IN2(n40), .IN3(n471), .IN4(n183), .IN5(n8), .IN6(n472), .QN(
          n469));
   OAI222X1 U878 (.IN1(n1546), .IN2(n36), .IN3(n475), .IN4(n331), .IN5(n1556), .IN6(n12), .
          QN(n474));
   NAND4X0 U879 (.IN1(n476), .IN2(n320), .IN3(n477), .IN4(n478), .QN(n473));
   AOI21X1 U880 (.IN1(n1569), .IN2(n391), .IN3(n355), .QN(n471));
   OA221X1 U881 (.IN1(n1552), .IN2(n1570), .IN3(n1569), .IN4(n1542), .IN5(n479), .Q(n470)
          );
   NAND4X0 U882 (.IN1(n481), .IN2(n478), .IN3(n482), .IN4(n483), .QN(n468));
   OA222X1 U883 (.IN1(n331), .IN2(n1558), .IN3(n39), .IN4(n475), .IN5(n1568), .IN6(n1556)
          , .Q(n483));
   NAND3X0 U884 (.IN1(n16), .IN2(n1568), .IN3(n340), .QN(n482));
   NAND3X0 U885 (.IN1(n390), .IN2(n484), .IN3(n485), .QN(n467));
   OA221X1 U886 (.IN1(n1570), .IN2(n1560), .IN3(n1568), .IN4(n1546), .IN5(n486), .Q(n485)
          );
   NAND3X0 U887 (.IN1(n342), .IN2(n1566), .IN3(n340), .QN(n486));
   OA22X1 U888 (.IN1(n1558), .IN2(n396), .IN3(n1542), .IN4(n1570), .Q(n390));
   AO221X1 U889 (.IN1(n373), .IN2(n487), .IN3(sboxw[6]), .IN4(n488), .IN5(n489), .Q(n465)
          );
   NAND4X0 U891 (.IN1(n491), .IN2(n321), .IN3(n492), .IN4(n493), .QN(n490));
   OA222X1 U892 (.IN1(n331), .IN2(n1556), .IN3(n1569), .IN4(n398), .IN5(n1570), .IN6(n1549)
          , .Q(n493));
   NAND3X0 U893 (.IN1(n1548), .IN2(n1568), .IN3(n16), .QN(n492));
   AO222X1 U894 (.IN1(n494), .IN2(n40), .IN3(n366), .IN4(n495), .IN5(n8), .IN6(n496), .Q(
          n488));
   NAND4X0 U895 (.IN1(n1542), .IN2(n393), .IN3(n497), .IN4(n498), .QN(n496));
   OA222X1 U896 (.IN1(n1547), .IN2(n1569), .IN3(n1568), .IN4(n499), .IN5(n1571), .IN6(
          n1560), .Q(n498));
   AO21X1 U897 (.IN1(n1552), .IN2(n397), .IN3(n35), .Q(n497));
   NAND3X0 U898 (.IN1(n500), .IN2(n1561), .IN3(n501), .QN(n495));
   NAND3X0 U899 (.IN1(n477), .IN2(n1550), .IN3(n502), .QN(n494));
   NAND4X0 U900 (.IN1(n328), .IN2(n1558), .IN3(n503), .IN4(n504), .QN(n487));
   OA22X1 U901 (.IN1(n7), .IN2(n1561), .IN3(n35), .IN4(n1557), .Q(n504));
   OR2X1 U902 (.IN1(n397), .IN2(n39), .Q(n503));
   AO221X1 U904 (.IN1(n309), .IN2(n508), .IN3(n307), .IN4(n509), .IN5(n510), .Q(n507));
   AO22X1 U905 (.IN1(n375), .IN2(n511), .IN3(n373), .IN4(n512), .Q(n510));
   NAND3X0 U906 (.IN1(n513), .IN2(n454), .IN3(n514), .QN(n512));
   OA22X1 U907 (.IN1(n1571), .IN2(n1555), .IN3(n1551), .IN4(n1569), .Q(n514));
   NAND3X0 U908 (.IN1(n370), .IN2(n1553), .IN3(n1563), .QN(n513));
   NAND4X0 U909 (.IN1(n515), .IN2(n423), .IN3(n516), .IN4(n517), .QN(n511));
   AOI222X1 U910 (.IN1(n447), .IN2(n417), .IN3(n1571), .IN4(n433), .IN5(n518), .IN6(n331)
          , .QN(n517));
   OA22X1 U911 (.IN1(n1566), .IN2(n39), .IN3(n1570), .IN4(n16), .Q(n417));
   OA22X1 U912 (.IN1(n1571), .IN2(n1556), .IN3(n1), .IN4(n1560), .Q(n516));
   NAND4X0 U913 (.IN1(n481), .IN2(n1552), .IN3(n422), .IN4(n519), .QN(n509));
   OA222X1 U914 (.IN1(n1563), .IN2(n1570), .IN3(n15), .IN4(n480), .IN5(n370), .IN6(n1556)
          , .Q(n519));
   NAND3X0 U915 (.IN1(n17), .IN2(n1566), .IN3(n35), .QN(n481));
   NAND4X0 U916 (.IN1(n352), .IN2(n491), .IN3(n521), .IN4(n522), .QN(n508));
   OA222X1 U917 (.IN1(n388), .IN2(n1552), .IN3(n1571), .IN4(n1560), .IN5(n1567), .IN6(
          n1545), .Q(n522));
   NAND3X0 U918 (.IN1(n1569), .IN2(n1553), .IN3(n1563), .QN(n521));
   NAND4X0 U919 (.IN1(n523), .IN2(n524), .IN3(n525), .IN4(n526), .QN(n506));
   OA222X1 U920 (.IN1(n527), .IN2(n40), .IN3(n8), .IN4(n528), .IN5(n1567), .IN6(n564), .Q(
          n526));
   NOR4X0 U921 (.IN1(n529), .IN2(n530), .IN3(n531), .IN4(n532), .QN(n527));
   AO222X1 U922 (.IN1(n518), .IN2(n1569), .IN3(n433), .IN4(n35), .IN5(n388), .IN6(n447), .
          Q(n529));
   OA22X1 U923 (.IN1(n15), .IN2(n16), .IN3(n1570), .IN4(n1566), .Q(n388));
   NAND3X0 U924 (.IN1(sboxw[1]), .IN2(n1548), .IN3(n366), .QN(n525));
   NAND3X0 U925 (.IN1(n15), .IN2(n17), .IN3(n327), .QN(n523));
   NAND4X0 U926 (.IN1(n524), .IN2(n454), .IN3(n533), .IN4(n534), .QN(n505));
   OA222X1 U927 (.IN1(n535), .IN2(n40), .IN3(n1561), .IN4(n325), .IN5(n39), .IN6(n564), .Q(
          n534));
   NOR4X0 U928 (.IN1(n536), .IN2(n537), .IN3(n538), .IN4(n539), .QN(n535));
   AO222X1 U929 (.IN1(n541), .IN2(n7), .IN3(n316), .IN4(n1569), .IN5(n386), .IN6(n1568), .
          Q(n536));
   NAND3X0 U930 (.IN1(n410), .IN2(n40), .IN3(n391), .QN(n524));
   AO222X1 U932 (.IN1(n548), .IN2(n549), .IN3(n550), .IN4(n551), .IN5(n552), .IN6(n49), .Q(
          n547));
   NAND4X0 U933 (.IN1(n553), .IN2(n554), .IN3(n555), .IN4(n556), .QN(n552));
   AOI222X1 U934 (.IN1(n557), .IN2(n14), .IN3(n558), .IN4(n88), .IN5(n11), .IN6(n559), .QN(
          n556));
   NAND4X0 U935 (.IN1(n560), .IN2(n62), .IN3(n561), .IN4(n562), .QN(n559));
   OA22X1 U936 (.IN1(n33), .IN2(n565), .IN3(n71), .IN4(n566), .Q(n555));
   NAND3X0 U937 (.IN1(n86), .IN2(n83), .IN3(n568), .QN(n553));
   NAND4X0 U938 (.IN1(n84), .IN2(n569), .IN3(n570), .IN4(n571), .QN(n551));
   OA222X1 U939 (.IN1(n572), .IN2(n70), .IN3(n90), .IN4(n573), .IN5(n34), .IN6(n68), .Q(
          n571));
   AND2X1 U940 (.IN1(n75), .IN2(n574), .Q(n570));
   NAND4X0 U941 (.IN1(n576), .IN2(n577), .IN3(n578), .IN4(n579), .QN(n549));
   OA22X1 U942 (.IN1(n580), .IN2(n90), .IN3(n89), .IN4(n75), .Q(n579));
   NAND3X0 U943 (.IN1(n33), .IN2(n25), .IN3(n581), .QN(n578));
   NAND3X0 U944 (.IN1(n26), .IN2(n582), .IN3(n583), .QN(n576));
   NAND4X0 U945 (.IN1(n584), .IN2(n50), .IN3(n585), .IN4(n586), .QN(n546));
   OA222X1 U946 (.IN1(n53), .IN2(n587), .IN3(n588), .IN4(n47), .IN5(n583), .IN6(n54), .Q(
          n586));
   AND3X1 U947 (.IN1(n589), .IN2(n69), .IN3(n569), .Q(n588));
   OA22X1 U948 (.IN1(n591), .IN2(n57), .IN3(n11), .IN4(n592), .Q(n585));
   AND3X1 U949 (.IN1(n593), .IN2(n594), .IN3(n595), .Q(n592));
   NOR3X0 U950 (.IN1(n596), .IN2(n597), .IN3(n598), .QN(n591));
   OA221X1 U951 (.IN1(n70), .IN2(n566), .IN3(n26), .IN4(n603), .IN5(n604), .Q(n602));
   OA22X1 U952 (.IN1(n572), .IN2(n59), .IN3(n57), .IN4(n88), .Q(n603));
   AOI222X1 U953 (.IN1(n11), .IN2(n605), .IN3(n606), .IN4(n47), .IN5(n596), .IN6(n607), .
          QN(n601));
   NAND3X0 U954 (.IN1(n608), .IN2(n609), .IN3(n610), .QN(n605));
   OA222X1 U955 (.IN1(n611), .IN2(n79), .IN3(n34), .IN4(n573), .IN5(n89), .IN6(n68), .Q(
          n610));
   AO222X1 U957 (.IN1(n614), .IN2(n615), .IN3(n616), .IN4(n617), .IN5(sboxw[30]), .IN6(
          n618), .Q(n613));
   AO221X1 U958 (.IN1(n11), .IN2(n619), .IN3(n620), .IN4(n47), .IN5(n621), .Q(n618));
   AO22X1 U959 (.IN1(n572), .IN2(n622), .IN3(n558), .IN4(n34), .Q(n621));
   OA221X1 U960 (.IN1(n583), .IN2(n65), .IN3(n24), .IN4(n625), .IN5(n626), .Q(n624));
   NAND3X0 U961 (.IN1(n85), .IN2(n72), .IN3(n611), .QN(n626));
   OA222X1 U962 (.IN1(n629), .IN2(n71), .IN3(n74), .IN4(n2), .IN5(n80), .IN6(n88), .Q(n623)
          );
   NAND3X0 U963 (.IN1(n630), .IN2(n594), .IN3(n631), .QN(n619));
   NAND4X0 U964 (.IN1(n633), .IN2(n634), .IN3(n635), .IN4(n636), .QN(n617));
   OA222X1 U965 (.IN1(n14), .IN2(n68), .IN3(n637), .IN4(n638), .IN5(n46), .IN6(n65), .Q(
          n636));
   OR2X1 U966 (.IN1(n639), .IN2(n24), .Q(n635));
   NAND4X0 U967 (.IN1(n574), .IN2(n68), .IN3(n640), .IN4(n641), .QN(n615));
   OA222X1 U968 (.IN1(sboxw[25]), .IN2(n71), .IN3(n86), .IN4(n64), .IN5(n583), .IN6(n74), .
          Q(n641));
   OA22X1 U969 (.IN1(n632), .IN2(n642), .IN3(n88), .IN4(n75), .Q(n640));
   AO221X1 U970 (.IN1(n548), .IN2(n643), .IN3(n644), .IN4(n49), .IN5(n645), .Q(n612));
   AO22X1 U971 (.IN1(n646), .IN2(sboxw[30]), .IN3(n550), .IN4(n647), .Q(n645));
   OA221X1 U972 (.IN1(n24), .IN2(n65), .IN3(n2), .IN4(n61), .IN5(n650), .Q(n649));
   AOI222X1 U973 (.IN1(n72), .IN2(n651), .IN3(n46), .IN4(n563), .IN5(n652), .IN6(n637), .
          QN(n648));
   OA221X1 U974 (.IN1(n655), .IN2(n53), .IN3(n656), .IN4(n59), .IN5(n78), .Q(n654));
   AND2X1 U975 (.IN1(n62), .IN2(n657), .Q(n655));
   OA222X1 U976 (.IN1(n658), .IN2(n76), .IN3(n659), .IN4(n47), .IN5(n11), .IN6(n660), .Q(
          n653));
   OA22X1 U977 (.IN1(n658), .IN2(n71), .IN3(sboxw[27]), .IN4(n611), .Q(n660));
   NAND4X0 U978 (.IN1(n661), .IN2(n662), .IN3(n663), .IN4(n664), .QN(n643));
   OR2X1 U979 (.IN1(n80), .IN2(n629), .Q(n662));
   AO221X1 U981 (.IN1(n375), .IN2(n668), .IN3(n309), .IN4(n669), .IN5(n670), .Q(n667));
   AO22X1 U982 (.IN1(n307), .IN2(n671), .IN3(n373), .IN4(n672), .Q(n670));
   NAND4X0 U983 (.IN1(n392), .IN2(n409), .IN3(n673), .IN4(n674), .QN(n672));
   OA222X1 U984 (.IN1(n396), .IN2(n1557), .IN3(sboxw[1]), .IN4(n1546), .IN5(n36), .IN6(
          n1560), .Q(n674));
   OA22X1 U985 (.IN1(n1567), .IN2(n499), .IN3(n1566), .IN4(n416), .Q(n673));
   NAND4X0 U986 (.IN1(n409), .IN2(n491), .IN3(n333), .IN4(n675), .QN(n671));
   OA22X1 U987 (.IN1(n1568), .IN2(n676), .IN3(n1570), .IN4(n499), .Q(n675));
   OA221X1 U988 (.IN1(sboxw[1]), .IN2(n1549), .IN3(n679), .IN4(n1570), .IN5(n680), .Q(n678)
          );
   OA222X1 U989 (.IN1(n1547), .IN2(n1), .IN3(n7), .IN4(n1560), .IN5(n1567), .IN6(n1558), .
          Q(n677));
   NAND4X0 U990 (.IN1(n491), .IN2(n478), .IN3(n681), .IN4(n682), .QN(n668));
   OA221X1 U991 (.IN1(sboxw[1]), .IN2(n1551), .IN3(n1567), .IN4(n1556), .IN5(n683), .Q(
          n682));
   AO221X1 U992 (.IN1(n684), .IN2(n39), .IN3(n8), .IN4(n685), .IN5(n686), .Q(n666));
   NAND3X0 U993 (.IN1(n1541), .IN2(n687), .IN3(n688), .QN(n686));
   NAND4X0 U995 (.IN1(n689), .IN2(n1559), .IN3(n690), .IN4(n691), .QN(n685));
   NAND3X0 U996 (.IN1(n341), .IN2(n1), .IN3(n17), .QN(n689));
   AO221X1 U997 (.IN1(n8), .IN2(n692), .IN3(n693), .IN4(n40), .IN5(n694), .Q(n665));
   AO221X1 U998 (.IN1(n359), .IN2(n1567), .IN3(n317), .IN4(n342), .IN5(n358), .Q(n694));
   NAND4X0 U999 (.IN1(n321), .IN2(n1555), .IN3(n695), .IN4(n696), .QN(n693));
   OA222X1 U1000 (.IN1(n1567), .IN2(n1549), .IN3(n697), .IN4(n39), .IN5(n1570), .IN6(n480)
          , .Q(n696));
   NAND3X0 U1001 (.IN1(n698), .IN2(n409), .IN3(n683), .QN(n692));
   OA22X1 U1002 (.IN1(n1555), .IN2(n39), .IN3(n1558), .IN4(n396), .Q(n683));
   AO222X1 U1003 (.IN1(n545), .IN2(n699), .IN3(n700), .IN4(n48), .IN5(n543), .IN6(n701), .
          Q(new_sboxw[29]));
   AO222X1 U1004 (.IN1(n607), .IN2(n702), .IN3(n703), .IN4(n47), .IN5(n11), .IN6(n704), .Q(
          n701));
   NAND4X0 U1005 (.IN1(n587), .IN2(n562), .IN3(n569), .IN4(n705), .QN(n704));
   OA221X1 U1006 (.IN1(n2), .IN2(n79), .IN3(n706), .IN4(n87), .IN5(n81), .Q(n705));
   NAND3X0 U1007 (.IN1(n63), .IN2(n561), .IN3(n709), .QN(n703));
   AO221X1 U1008 (.IN1(n26), .IN2(n87), .IN3(n90), .IN4(n72), .IN5(n83), .Q(n702));
   AO22X1 U1009 (.IN1(n710), .IN2(n49), .IN3(sboxw[30]), .IN4(n711), .Q(n700));
   AO221X1 U1010 (.IN1(n607), .IN2(n712), .IN3(n11), .IN4(n713), .IN5(n714), .Q(n711));
   AO22X1 U1011 (.IN1(n715), .IN2(n24), .IN3(n716), .IN4(n568), .Q(n714));
   NAND4X0 U1012 (.IN1(n594), .IN2(n717), .IN3(n718), .IN4(n719), .QN(n713));
   OA221X1 U1013 (.IN1(n46), .IN2(n75), .IN3(n637), .IN4(n68), .IN5(n720), .Q(n719));
   AO222X1 U1014 (.IN1(n637), .IN2(n632), .IN3(n33), .IN4(n722), .IN5(n652), .IN6(n89), .Q(
          n712));
   NAND4X0 U1015 (.IN1(n73), .IN2(n717), .IN3(n723), .IN4(n724), .QN(n710));
   OA221X1 U1016 (.IN1(n725), .IN2(n47), .IN3(n11), .IN4(n726), .IN5(n727), .Q(n724));
   OA22X1 U1017 (.IN1(n728), .IN2(n53), .IN3(n637), .IN4(n75), .Q(n727));
   AND3X1 U1018 (.IN1(n63), .IN2(n80), .IN3(n657), .Q(n728));
   NAND4X0 U1019 (.IN1(n554), .IN2(n577), .IN3(n731), .IN4(n732), .QN(n699));
   OA222X1 U1020 (.IN1(n733), .IN2(n47), .IN3(n11), .IN4(n734), .IN5(n54), .IN6(n2), .Q(
          n732));
   OA22X1 U1021 (.IN1(n64), .IN2(sboxw[25]), .IN3(n77), .IN4(n583), .Q(n608));
   OA221X1 U1022 (.IN1(n46), .IN2(n80), .IN3(n34), .IN4(n70), .IN5(n736), .Q(n733));
   OA22X1 U1023 (.IN1(n53), .IN2(n737), .IN3(n738), .IN4(n57), .Q(n731));
   NAND3X0 U1024 (.IN1(n739), .IN2(n2), .IN3(n632), .QN(n554));
   AO222X1 U1026 (.IN1(n614), .IN2(n742), .IN3(n616), .IN4(n743), .IN5(sboxw[30]), .IN6(
          n744), .Q(n741));
   OAI222X1 U1027 (.IN1(n745), .IN2(n47), .IN3(n746), .IN4(n53), .IN5(n11), .IN6(n747), .
          QN(n744));
   OAI222X1 U1028 (.IN1(n65), .IN2(n34), .IN3(n750), .IN4(n572), .IN5(n75), .IN6(n14), .QN(
          n749));
   NAND4X0 U1029 (.IN1(n751), .IN2(n561), .IN3(n752), .IN4(n753), .QN(n748));
   AOI21X1 U1030 (.IN1(n88), .IN2(n632), .IN3(n596), .QN(n746));
   OA221X1 U1031 (.IN1(n71), .IN2(n89), .IN3(n88), .IN4(n61), .IN5(n754), .Q(n745));
   NAND4X0 U1032 (.IN1(n756), .IN2(n753), .IN3(n757), .IN4(n758), .QN(n743));
   OA222X1 U1033 (.IN1(n572), .IN2(n77), .IN3(n46), .IN4(n750), .IN5(n87), .IN6(n75), .Q(
          n758));
   NAND3X0 U1034 (.IN1(n25), .IN2(n87), .IN3(n581), .QN(n757));
   NAND3X0 U1035 (.IN1(n631), .IN2(n759), .IN3(n760), .QN(n742));
   OA221X1 U1036 (.IN1(n89), .IN2(n79), .IN3(n87), .IN4(n65), .IN5(n761), .Q(n760));
   NAND3X0 U1037 (.IN1(n5), .IN2(n85), .IN3(n581), .QN(n761));
   OA22X1 U1038 (.IN1(n77), .IN2(n637), .IN3(n61), .IN4(n89), .Q(n631));
   AO221X1 U1039 (.IN1(n614), .IN2(n762), .IN3(sboxw[30]), .IN4(n763), .IN5(n764), .Q(n740)
          );
   AO22X1 U1040 (.IN1(n616), .IN2(n765), .IN3(n611), .IN4(n622), .Q(n764));
   NAND4X0 U1041 (.IN1(n766), .IN2(n562), .IN3(n767), .IN4(n768), .QN(n765));
   OA222X1 U1042 (.IN1(n572), .IN2(n75), .IN3(n88), .IN4(n639), .IN5(n89), .IN6(n68), .Q(
          n768));
   NAND3X0 U1043 (.IN1(n67), .IN2(n87), .IN3(n25), .QN(n767));
   AO222X1 U1044 (.IN1(n769), .IN2(n47), .IN3(n607), .IN4(n770), .IN5(n11), .IN6(n771), .Q(
          n763));
   NAND4X0 U1045 (.IN1(n61), .IN2(n634), .IN3(n772), .IN4(n773), .QN(n771));
   OA222X1 U1046 (.IN1(n66), .IN2(n88), .IN3(n87), .IN4(n774), .IN5(n90), .IN6(n79), .Q(
          n773));
   AO21X1 U1047 (.IN1(n71), .IN2(n638), .IN3(n33), .Q(n772));
   NAND3X0 U1048 (.IN1(n775), .IN2(n80), .IN3(n776), .QN(n770));
   NAND3X0 U1049 (.IN1(n752), .IN2(n69), .IN3(n777), .QN(n769));
   NAND4X0 U1050 (.IN1(n569), .IN2(n77), .IN3(n778), .IN4(n779), .QN(n762));
   OA22X1 U1051 (.IN1(n5), .IN2(n80), .IN3(n33), .IN4(n76), .Q(n779));
   OR2X1 U1052 (.IN1(n638), .IN2(n46), .Q(n778));
   AO222X1 U1053 (.IN1(n543), .IN2(n780), .IN3(n545), .IN4(n781), .IN5(n782), .IN6(n48), .
          Q(new_sboxw[27]));
   AO221X1 U1054 (.IN1(n550), .IN2(n783), .IN3(n548), .IN4(n784), .IN5(n785), .Q(n782));
   AO22X1 U1055 (.IN1(n616), .IN2(n786), .IN3(n614), .IN4(n787), .Q(n785));
   NAND3X0 U1056 (.IN1(n788), .IN2(n729), .IN3(n789), .QN(n787));
   OA22X1 U1057 (.IN1(n90), .IN2(n74), .IN3(n70), .IN4(n88), .Q(n789));
   NAND3X0 U1058 (.IN1(n611), .IN2(n72), .IN3(n82), .QN(n788));
   NAND4X0 U1059 (.IN1(n790), .IN2(n664), .IN3(n791), .IN4(n792), .QN(n786));
   AOI222X1 U1060 (.IN1(n722), .IN2(n658), .IN3(n90), .IN4(n708), .IN5(n793), .IN6(n572), .
          QN(n792));
   OA22X1 U1061 (.IN1(n85), .IN2(n46), .IN3(n89), .IN4(n25), .Q(n658));
   OA22X1 U1062 (.IN1(n90), .IN2(n75), .IN3(n2), .IN4(n79), .Q(n791));
   NAND4X0 U1063 (.IN1(n756), .IN2(n71), .IN3(n663), .IN4(n794), .QN(n784));
   OA222X1 U1064 (.IN1(n82), .IN2(n89), .IN3(n24), .IN4(n755), .IN5(n611), .IN6(n75), .Q(
          n794));
   NAND3X0 U1065 (.IN1(n26), .IN2(n85), .IN3(n33), .QN(n756));
   NAND4X0 U1066 (.IN1(n593), .IN2(n766), .IN3(n796), .IN4(n797), .QN(n783));
   OA222X1 U1067 (.IN1(n629), .IN2(n71), .IN3(n90), .IN4(n79), .IN5(n86), .IN6(n64), .Q(
          n797));
   NAND3X0 U1068 (.IN1(n88), .IN2(n72), .IN3(n82), .QN(n796));
   NAND4X0 U1069 (.IN1(n798), .IN2(n799), .IN3(n800), .IN4(n801), .QN(n781));
   OA222X1 U1070 (.IN1(n802), .IN2(n47), .IN3(n11), .IN4(n803), .IN5(n86), .IN6(n58), .Q(
          n801));
   NOR4X0 U1071 (.IN1(n804), .IN2(n805), .IN3(n806), .IN4(n807), .QN(n802));
   AO222X1 U1072 (.IN1(n793), .IN2(n88), .IN3(n708), .IN4(n33), .IN5(n629), .IN6(n722), .Q(
          n804));
   OA22X1 U1073 (.IN1(n24), .IN2(n25), .IN3(n89), .IN4(n85), .Q(n629));
   NAND3X0 U1074 (.IN1(sboxw[25]), .IN2(n67), .IN3(n607), .QN(n800));
   NAND3X0 U1075 (.IN1(n24), .IN2(n26), .IN3(n568), .QN(n798));
   NAND4X0 U1076 (.IN1(n799), .IN2(n729), .IN3(n808), .IN4(n809), .QN(n780));
   OA222X1 U1077 (.IN1(n810), .IN2(n47), .IN3(n80), .IN4(n566), .IN5(n46), .IN6(n58), .Q(
          n809));
   NOR4X0 U1078 (.IN1(n811), .IN2(n812), .IN3(n813), .IN4(n814), .QN(n810));
   AO222X1 U1079 (.IN1(n816), .IN2(n5), .IN3(n557), .IN4(n88), .IN5(n627), .IN6(n87), .Q(
          n811));
   NAND3X0 U1080 (.IN1(n651), .IN2(n47), .IN3(n632), .QN(n799));
   AO222X1 U1081 (.IN1(n543), .IN2(n818), .IN3(n545), .IN4(n819), .IN5(n820), .IN6(n48), .
          Q(new_sboxw[26]));
   AO221X1 U1082 (.IN1(n616), .IN2(n821), .IN3(n550), .IN4(n822), .IN5(n823), .Q(n820));
   AO22X1 U1083 (.IN1(n548), .IN2(n824), .IN3(n614), .IN4(n825), .Q(n823));
   NAND4X0 U1084 (.IN1(n633), .IN2(n650), .IN3(n826), .IN4(n827), .QN(n825));
   OA222X1 U1085 (.IN1(n637), .IN2(n76), .IN3(sboxw[25]), .IN4(n65), .IN5(n34), .IN6(n79)
          , .Q(n827));
   OA22X1 U1086 (.IN1(n86), .IN2(n774), .IN3(n85), .IN4(n657), .Q(n826));
   NAND4X0 U1087 (.IN1(n650), .IN2(n766), .IN3(n574), .IN4(n828), .QN(n824));
   OA22X1 U1088 (.IN1(n87), .IN2(n829), .IN3(n89), .IN4(n774), .Q(n828));
   OA221X1 U1089 (.IN1(sboxw[25]), .IN2(n68), .IN3(n832), .IN4(n89), .IN5(n833), .Q(n831)
          );
   OA222X1 U1090 (.IN1(n66), .IN2(n2), .IN3(n583), .IN4(n79), .IN5(n86), .IN6(n77), .Q(
          n830));
   NAND4X0 U1091 (.IN1(n766), .IN2(n753), .IN3(n834), .IN4(n835), .QN(n821));
   OA221X1 U1092 (.IN1(sboxw[25]), .IN2(n70), .IN3(n86), .IN4(n75), .IN5(n836), .Q(n835)
          );
   AO221X1 U1093 (.IN1(n837), .IN2(n46), .IN3(n11), .IN4(n838), .IN5(n839), .Q(n819));
   NAND3X0 U1094 (.IN1(n60), .IN2(n840), .IN3(n841), .QN(n839));
   NAND3X0 U1095 (.IN1(n87), .IN2(n66), .IN3(n607), .QN(n841));
   NAND4X0 U1096 (.IN1(n842), .IN2(n78), .IN3(n843), .IN4(n844), .QN(n838));
   NAND3X0 U1097 (.IN1(n582), .IN2(n2), .IN3(n26), .QN(n842));
   AO221X1 U1098 (.IN1(n11), .IN2(n845), .IN3(n846), .IN4(n47), .IN5(n847), .Q(n818));
   AO221X1 U1099 (.IN1(n600), .IN2(n86), .IN3(n558), .IN4(n5), .IN5(n599), .Q(n847));
   NAND4X0 U1100 (.IN1(n562), .IN2(n74), .IN3(n848), .IN4(n849), .QN(n846));
   OA222X1 U1101 (.IN1(n86), .IN2(n68), .IN3(n850), .IN4(n46), .IN5(n89), .IN6(n755), .Q(
          n849));
   NAND3X0 U1102 (.IN1(n851), .IN2(n650), .IN3(n836), .QN(n845));
   OA22X1 U1103 (.IN1(n74), .IN2(n46), .IN3(n77), .IN4(n637), .Q(n836));
   AO222X1 U1105 (.IN1(n548), .IN2(n854), .IN3(n550), .IN4(n855), .IN5(n856), .IN6(n49), .
          Q(n853));
   NAND4X0 U1106 (.IN1(n857), .IN2(n567), .IN3(n858), .IN4(n859), .QN(n856));
   OA221X1 U1107 (.IN1(n575), .IN2(n76), .IN3(n776), .IN4(n57), .IN5(n860), .Q(n859));
   OA22X1 U1108 (.IN1(n637), .IN2(n51), .IN3(n87), .IN4(n58), .Q(n860));
   OA22X1 U1109 (.IN1(n46), .IN2(n83), .IN3(n66), .IN4(sboxw[25]), .Q(n776));
   OA22X1 U1110 (.IN1(n85), .IN2(n33), .IN3(n611), .IN4(n25), .Q(n575));
   OA22X1 U1111 (.IN1(n861), .IN2(n47), .IN3(n572), .IN4(n52), .Q(n858));
   OA22X1 U1112 (.IN1(n90), .IN2(n64), .IN3(n34), .IN4(n70), .Q(n861));
   NAND3X0 U1113 (.IN1(n90), .IN2(n47), .IN3(n628), .QN(n857));
   NAND4X0 U1114 (.IN1(n752), .IN2(n577), .IN3(n862), .IN4(n863), .QN(n855));
   OA222X1 U1115 (.IN1(n64), .IN2(n88), .IN3(n86), .IN4(n68), .IN5(n87), .IN6(n77), .Q(
          n863));
   OA22X1 U1116 (.IN1(n572), .IN2(n832), .IN3(n90), .IN4(n65), .Q(n862));
   NAND4X0 U1117 (.IN1(n73), .IN2(n595), .IN3(n864), .IN4(n865), .QN(n854));
   OA222X1 U1118 (.IN1(n86), .IN2(n80), .IN3(n88), .IN4(n65), .IN5(n64), .IN6(n2), .Q(n865)
          );
   OA22X1 U1119 (.IN1(n90), .IN2(n866), .IN3(n34), .IN4(n750), .Q(n864));
   AO221X1 U1120 (.IN1(n548), .IN2(n867), .IN3(n868), .IN4(n49), .IN5(n869), .Q(n852));
   AO22X1 U1121 (.IN1(n550), .IN2(n870), .IN3(n871), .IN4(n558), .Q(n869));
   NAND4X0 U1122 (.IN1(n720), .IN2(n751), .IN3(n872), .IN4(n873), .QN(n870));
   OA22X1 U1123 (.IN1(n33), .IN2(n64), .IN3(n71), .IN4(n2), .Q(n873));
   AO222X1 U1124 (.IN1(n739), .IN2(n874), .IN3(n11), .IN4(n875), .IN5(n876), .IN6(n47), .Q(
          n868));
   NAND3X0 U1125 (.IN1(n877), .IN2(n661), .IN3(n878), .QN(n876));
   OA222X1 U1126 (.IN1(n85), .IN2(n657), .IN3(n87), .IN4(n573), .IN5(sboxw[25]), .IN6(n61)
          , .Q(n878));
   OA22X1 U1127 (.IN1(n86), .IN2(n79), .IN3(n637), .IN4(n74), .Q(n877));
   NAND3X0 U1128 (.IN1(n717), .IN2(n753), .IN3(n593), .QN(n875));
   AO221X1 U1129 (.IN1(n632), .IN2(n88), .IN3(n24), .IN4(n652), .IN5(n879), .Q(n874));
   AO22X1 U1130 (.IN1(n590), .IN2(n87), .IN3(n722), .IN4(n90), .Q(n879));
   OA222X1 U1131 (.IN1(n87), .IN2(n68), .IN3(n882), .IN4(n90), .IN5(n583), .IN6(n832), .Q(
          n881));
   OA222X1 U1132 (.IN1(n80), .IN2(n2), .IN3(n24), .IN4(n77), .IN5(n572), .IN6(n64), .Q(
          n880));
   AO22X1 U1133 (.IN1(sboxw[31]), .IN2(n883), .IN3(n884), .IN4(n48), .Q(new_sboxw[24]));
   AO22X1 U1134 (.IN1(n885), .IN2(n49), .IN3(sboxw[30]), .IN4(n886), .Q(n884));
   NAND4X0 U1135 (.IN1(n887), .IN2(n55), .IN3(n888), .IN4(n889), .QN(n886));
   AOI222X1 U1136 (.IN1(n11), .IN2(n890), .IN3(n891), .IN4(n47), .IN5(n735), .IN6(n46), .
          QN(n889));
   NAND3X0 U1137 (.IN1(n587), .IN2(n594), .IN3(n892), .QN(n891));
   NAND4X0 U1138 (.IN1(n717), .IN2(n74), .IN3(n894), .IN4(n895), .QN(n890));
   OA222X1 U1139 (.IN1(n90), .IN2(n76), .IN3(n87), .IN4(n755), .IN5(n2), .IN6(n68), .Q(
          n895));
   OR2X1 U1140 (.IN1(n774), .IN2(n90), .Q(n833));
   NAND3X0 U1141 (.IN1(n33), .IN2(n26), .IN3(n568), .QN(n887));
   NAND4X0 U1142 (.IN1(n897), .IN2(n840), .IN3(n898), .IN4(n899), .QN(n885));
   AOI222X1 U1143 (.IN1(n11), .IN2(n900), .IN3(n715), .IN4(n88), .IN5(n735), .IN6(n89), .
          QN(n899));
   NAND4X0 U1144 (.IN1(n848), .IN2(n753), .IN3(n901), .IN4(n902), .QN(n900));
   OA222X1 U1145 (.IN1(n637), .IN2(n70), .IN3(n34), .IN4(n75), .IN5(n611), .IN6(n77), .Q(
          n902));
   NAND3X0 U1146 (.IN1(n88), .IN2(n85), .IN3(n67), .QN(n848));
   NAND3X0 U1147 (.IN1(n583), .IN2(n67), .IN3(n568), .QN(n897));
   AO222X1 U1148 (.IN1(sboxw[30]), .IN2(n903), .IN3(n548), .IN4(n904), .IN5(n905), .IN6(
          n49), .Q(n883));
   AO221X1 U1149 (.IN1(n906), .IN2(n47), .IN3(n627), .IN4(n611), .IN5(n907), .Q(n905));
   AO222X1 U1150 (.IN1(n600), .IN2(n89), .IN3(n908), .IN4(n25), .IN5(n607), .IN6(n909), .Q(
          n907));
   AO221X1 U1151 (.IN1(n583), .IN2(n722), .IN3(n632), .IN4(n90), .IN5(n721), .Q(n909));
   OAI221X1 U1152 (.IN1(n77), .IN2(n572), .IN3(n74), .IN4(n637), .IN5(n751), .QN(n906));
   AO221X1 U1153 (.IN1(n611), .IN2(n628), .IN3(n590), .IN4(n893), .IN5(n597), .Q(n904));
   XNOR2X1 U1154 (.IN1(n25), .IN2(n24), .Q(n911));
   AO221X1 U1155 (.IN1(n912), .IN2(n637), .IN3(n11), .IN4(n913), .IN5(n817), .Q(n903));
   NAND4X0 U1156 (.IN1(n69), .IN2(n68), .IN3(n914), .IN4(n915), .QN(n913));
   OA221X1 U1157 (.IN1(n14), .IN2(n74), .IN3(n64), .IN4(n88), .IN5(n916), .Q(n915));
   OA22X1 U1158 (.IN1(n611), .IN2(n79), .IN3(n90), .IN4(n77), .Q(n916));
   AO222X1 U1159 (.IN1(n917), .IN2(n918), .IN3(n919), .IN4(n920), .IN5(n921), .IN6(n91), .
          Q(new_sboxw[23]));
   AO222X1 U1160 (.IN1(n922), .IN2(n923), .IN3(n924), .IN4(n925), .IN5(n926), .IN6(n92), .
          Q(n921));
   NAND4X0 U1161 (.IN1(n927), .IN2(n928), .IN3(n929), .IN4(n930), .QN(n926));
   AOI222X1 U1162 (.IN1(n931), .IN2(n13), .IN3(n932), .IN4(n131), .IN5(n10), .IN6(n933), .
          QN(n930));
   NAND4X0 U1163 (.IN1(n934), .IN2(n105), .IN3(n935), .IN4(n936), .QN(n933));
   OA22X1 U1164 (.IN1(n31), .IN2(n939), .IN3(n114), .IN4(n940), .Q(n929));
   NAND4X0 U1166 (.IN1(n127), .IN2(n943), .IN3(n944), .IN4(n945), .QN(n925));
   AND2X1 U1168 (.IN1(n118), .IN2(n948), .Q(n944));
   NAND4X0 U1169 (.IN1(n950), .IN2(n951), .IN3(n952), .IN4(n953), .QN(n923));
   OA22X1 U1170 (.IN1(n954), .IN2(n133), .IN3(n132), .IN4(n118), .Q(n953));
   NAND3X0 U1171 (.IN1(n31), .IN2(n22), .IN3(n955), .QN(n952));
   NAND4X0 U1173 (.IN1(n958), .IN2(n93), .IN3(n959), .IN4(n960), .QN(n920));
   OA222X1 U1174 (.IN1(n96), .IN2(n961), .IN3(n962), .IN4(n45), .IN5(n957), .IN6(n97), .Q(
          n960));
   AND3X1 U1175 (.IN1(n963), .IN2(n112), .IN3(n943), .Q(n962));
   OA22X1 U1176 (.IN1(n965), .IN2(n100), .IN3(n10), .IN4(n966), .Q(n959));
   AND3X1 U1177 (.IN1(n967), .IN2(n968), .IN3(n969), .Q(n966));
   NOR3X0 U1178 (.IN1(n970), .IN2(n971), .IN3(n972), .QN(n965));
   OA221X1 U1179 (.IN1(n113), .IN2(n940), .IN3(n23), .IN4(n977), .IN5(n978), .Q(n976));
   OA22X1 U1180 (.IN1(n946), .IN2(n102), .IN3(n100), .IN4(n131), .Q(n977));
   AOI222X1 U1181 (.IN1(n10), .IN2(n979), .IN3(n980), .IN4(n45), .IN5(n970), .IN6(n981), .
          QN(n975));
   NAND3X0 U1182 (.IN1(n982), .IN2(n983), .IN3(n984), .QN(n979));
   OA222X1 U1183 (.IN1(n985), .IN2(n122), .IN3(n31), .IN4(n947), .IN5(n132), .IN6(n111), .
          Q(n984));
   AO22X1 U1184 (.IN1(n986), .IN2(n91), .IN3(sboxw[23]), .IN4(n987), .Q(new_sboxw[22]));
   AO222X1 U1185 (.IN1(n988), .IN2(n989), .IN3(n990), .IN4(n991), .IN5(sboxw[22]), .IN6(
          n992), .Q(n987));
   AO221X1 U1186 (.IN1(n10), .IN2(n993), .IN3(n994), .IN4(n45), .IN5(n995), .Q(n992));
   AO22X1 U1187 (.IN1(n946), .IN2(n996), .IN3(n932), .IN4(n31), .Q(n995));
   NAND3X0 U1189 (.IN1(n128), .IN2(n115), .IN3(n985), .QN(n1000));
   OA222X1 U1190 (.IN1(n1003), .IN2(n114), .IN3(n117), .IN4(n32), .IN5(n123), .IN6(n131), .
          Q(n997));
   NAND3X0 U1191 (.IN1(n1004), .IN2(n968), .IN3(n1005), .QN(n993));
   NAND4X0 U1192 (.IN1(n1007), .IN2(n1008), .IN3(n1009), .IN4(n1010), .QN(n991));
   OA222X1 U1193 (.IN1(sboxw[17]), .IN2(n111), .IN3(n1011), .IN4(n1012), .IN5(n44), .IN6(
          n108), .Q(n1010));
   OR2X1 U1194 (.IN1(n1013), .IN2(n21), .Q(n1009));
   NAND4X0 U1195 (.IN1(n948), .IN2(n111), .IN3(n1014), .IN4(n1015), .QN(n989));
   OA222X1 U1196 (.IN1(sboxw[17]), .IN2(n114), .IN3(n129), .IN4(n107), .IN5(n957), .IN6(
          n117), .Q(n1015));
   OA22X1 U1197 (.IN1(n1006), .IN2(n1016), .IN3(n131), .IN4(n118), .Q(n1014));
   AO221X1 U1198 (.IN1(n922), .IN2(n1017), .IN3(n1018), .IN4(n92), .IN5(n1019), .Q(n986)
          );
   AO22X1 U1199 (.IN1(n1020), .IN2(sboxw[22]), .IN3(n924), .IN4(n1021), .Q(n1019));
   OA221X1 U1200 (.IN1(n21), .IN2(n108), .IN3(n32), .IN4(n104), .IN5(n1024), .Q(n1023));
   AOI222X1 U1201 (.IN1(n115), .IN2(n1025), .IN3(n44), .IN4(n937), .IN5(n1026), .IN6(n1011)
          , .QN(n1022));
   OA221X1 U1202 (.IN1(n1029), .IN2(n96), .IN3(n1030), .IN4(n102), .IN5(n121), .Q(n1028)
          );
   AND2X1 U1203 (.IN1(n105), .IN2(n1031), .Q(n1029));
   OA222X1 U1204 (.IN1(n1032), .IN2(n119), .IN3(n1033), .IN4(n45), .IN5(n10), .IN6(n1034)
          , .Q(n1027));
   OA22X1 U1205 (.IN1(n1032), .IN2(n114), .IN3(sboxw[19]), .IN4(n985), .Q(n1034));
   NAND4X0 U1206 (.IN1(n1035), .IN2(n1036), .IN3(n1037), .IN4(n1038), .QN(n1017));
   OR2X1 U1207 (.IN1(n123), .IN2(n1003), .Q(n1036));
   AO222X1 U1209 (.IN1(n981), .IN2(n1042), .IN3(n1043), .IN4(n45), .IN5(n10), .IN6(n1044)
          , .Q(n1041));
   NAND4X0 U1210 (.IN1(n961), .IN2(n936), .IN3(n943), .IN4(n1045), .QN(n1044));
   OA221X1 U1211 (.IN1(n32), .IN2(n122), .IN3(n1046), .IN4(n130), .IN5(n124), .Q(n1045));
   NAND3X0 U1212 (.IN1(n106), .IN2(n935), .IN3(n1049), .QN(n1043));
   AO221X1 U1213 (.IN1(n23), .IN2(n130), .IN3(n133), .IN4(n115), .IN5(n126), .Q(n1042));
   AO22X1 U1216 (.IN1(n1055), .IN2(n21), .IN3(n1056), .IN4(n942), .Q(n1054));
   NAND4X0 U1217 (.IN1(n968), .IN2(n1057), .IN3(n1058), .IN4(n1059), .QN(n1053));
   OA221X1 U1218 (.IN1(n44), .IN2(n118), .IN3(n1011), .IN4(n111), .IN5(n1060), .Q(n1059)
          );
   AO222X1 U1219 (.IN1(n1011), .IN2(n1006), .IN3(n31), .IN4(n1062), .IN5(n1026), .IN6(n132)
          , .Q(n1052));
   NAND4X0 U1220 (.IN1(n116), .IN2(n1057), .IN3(n1063), .IN4(n1064), .QN(n1050));
   OA221X1 U1221 (.IN1(n1065), .IN2(n45), .IN3(n10), .IN4(n1066), .IN5(n1067), .Q(n1064)
          );
   OA22X1 U1222 (.IN1(n1068), .IN2(n96), .IN3(n1011), .IN4(n118), .Q(n1067));
   AND3X1 U1223 (.IN1(n106), .IN2(n123), .IN3(n1031), .Q(n1068));
   NAND4X0 U1224 (.IN1(n928), .IN2(n951), .IN3(n1071), .IN4(n1072), .QN(n1039));
   OA222X1 U1225 (.IN1(n1073), .IN2(n45), .IN3(n10), .IN4(n1074), .IN5(n97), .IN6(n32), .Q(
          n1072));
   OA22X1 U1226 (.IN1(n107), .IN2(sboxw[17]), .IN3(n120), .IN4(n957), .Q(n982));
   OA221X1 U1227 (.IN1(n44), .IN2(n123), .IN3(n31), .IN4(n113), .IN5(n1076), .Q(n1073));
   OA22X1 U1228 (.IN1(n96), .IN2(n1077), .IN3(n1078), .IN4(n100), .Q(n1071));
   NAND3X0 U1229 (.IN1(n1079), .IN2(n32), .IN3(n1006), .QN(n928));
   AO22X1 U1230 (.IN1(n1080), .IN2(n91), .IN3(sboxw[23]), .IN4(n1081), .Q(new_sboxw[20])
          );
   AO222X1 U1231 (.IN1(n988), .IN2(n1082), .IN3(n990), .IN4(n1083), .IN5(sboxw[22]), .IN6(
          n1084), .Q(n1081));
   OAI222X1 U1232 (.IN1(n1085), .IN2(n45), .IN3(n1086), .IN4(n96), .IN5(n10), .IN6(n1087)
          , .QN(n1084));
   NAND4X0 U1234 (.IN1(n1091), .IN2(n935), .IN3(n1092), .IN4(n1093), .QN(n1088));
   AOI21X1 U1235 (.IN1(n131), .IN2(n1006), .IN3(n970), .QN(n1086));
   OA221X1 U1236 (.IN1(n114), .IN2(n132), .IN3(n131), .IN4(n104), .IN5(n1094), .Q(n1085)
          );
   NAND4X0 U1237 (.IN1(n1096), .IN2(n1093), .IN3(n1097), .IN4(n1098), .QN(n1083));
   OA222X1 U1238 (.IN1(n946), .IN2(n120), .IN3(n44), .IN4(n1090), .IN5(n130), .IN6(n118), .
          Q(n1098));
   NAND3X0 U1239 (.IN1(n22), .IN2(n130), .IN3(n955), .QN(n1097));
   NAND3X0 U1240 (.IN1(n1005), .IN2(n1099), .IN3(n1100), .QN(n1082));
   OA221X1 U1241 (.IN1(n132), .IN2(n122), .IN3(n130), .IN4(n108), .IN5(n1101), .Q(n1100)
          );
   OA22X1 U1243 (.IN1(n120), .IN2(n1011), .IN3(n104), .IN4(n132), .Q(n1005));
   NAND4X0 U1246 (.IN1(n1106), .IN2(n936), .IN3(n1107), .IN4(n1108), .QN(n1105));
   OA222X1 U1247 (.IN1(n946), .IN2(n118), .IN3(n131), .IN4(n1013), .IN5(n132), .IN6(n111)
          , .Q(n1108));
   NAND3X0 U1248 (.IN1(n110), .IN2(n130), .IN3(n22), .QN(n1107));
   AO222X1 U1249 (.IN1(n1109), .IN2(n45), .IN3(n981), .IN4(n1110), .IN5(n10), .IN6(n1111)
          , .Q(n1103));
   NAND4X0 U1250 (.IN1(n104), .IN2(n1008), .IN3(n1112), .IN4(n1113), .QN(n1111));
   OA222X1 U1251 (.IN1(n109), .IN2(n131), .IN3(n130), .IN4(n1114), .IN5(n133), .IN6(n122)
          , .Q(n1113));
   AO21X1 U1252 (.IN1(n114), .IN2(n1012), .IN3(n31), .Q(n1112));
   NAND3X0 U1253 (.IN1(n1115), .IN2(n123), .IN3(n1116), .QN(n1110));
   NAND3X0 U1254 (.IN1(n1092), .IN2(n112), .IN3(n1117), .QN(n1109));
   NAND4X0 U1255 (.IN1(n943), .IN2(n120), .IN3(n1118), .IN4(n1119), .QN(n1102));
   OA22X1 U1256 (.IN1(n957), .IN2(n123), .IN3(n938), .IN4(n119), .Q(n1119));
   OR2X1 U1257 (.IN1(n1012), .IN2(n44), .Q(n1118));
   AO222X1 U1259 (.IN1(n307), .IN2(n1122), .IN3(n309), .IN4(n1123), .IN5(n1124), .IN6(n179)
          , .Q(n1121));
   NAND4X0 U1260 (.IN1(n1125), .IN2(n326), .IN3(n1126), .IN4(n1127), .QN(n1124));
   OA221X1 U1261 (.IN1(n334), .IN2(n1557), .IN3(n501), .IN4(n323), .IN5(n1128), .Q(n1127)
          );
   OA22X1 U1262 (.IN1(n396), .IN2(n181), .IN3(n1568), .IN4(n564), .Q(n1128));
   OA22X1 U1263 (.IN1(n39), .IN2(n1564), .IN3(n1547), .IN4(sboxw[1]), .Q(n501));
   OA22X1 U1264 (.IN1(n1566), .IN2(n35), .IN3(n370), .IN4(n16), .Q(n334));
   OA22X1 U1265 (.IN1(n1129), .IN2(n40), .IN3(n331), .IN4(n182), .Q(n1126));
   OA22X1 U1266 (.IN1(n1571), .IN2(n1545), .IN3(n36), .IN4(n1551), .Q(n1129));
   NAND3X0 U1267 (.IN1(n1571), .IN2(n40), .IN3(n387), .QN(n1125));
   NAND4X0 U1268 (.IN1(n477), .IN2(n336), .IN3(n1130), .IN4(n1131), .QN(n1123));
   OA222X1 U1269 (.IN1(n1545), .IN2(n1569), .IN3(n1567), .IN4(n1549), .IN5(n1568), .IN6(
          n1558), .Q(n1131));
   OA22X1 U1270 (.IN1(n331), .IN2(n679), .IN3(n1571), .IN4(n1546), .Q(n1130));
   NAND4X0 U1271 (.IN1(n1554), .IN2(n354), .IN3(n1132), .IN4(n1133), .QN(n1122));
   OA222X1 U1272 (.IN1(n1567), .IN2(n1561), .IN3(n1569), .IN4(n1546), .IN5(n1545), .IN6(n1)
          , .Q(n1133));
   OA22X1 U1273 (.IN1(n1571), .IN2(n1134), .IN3(n36), .IN4(n475), .Q(n1132));
   AO221X1 U1274 (.IN1(n307), .IN2(n1135), .IN3(n1136), .IN4(n179), .IN5(n1137), .Q(n1120)
          );
   AO22X1 U1275 (.IN1(n309), .IN2(n1138), .IN3(n1139), .IN4(n317), .Q(n1137));
   NAND4X0 U1276 (.IN1(n445), .IN2(n476), .IN3(n1140), .IN4(n1141), .QN(n1138));
   OA22X1 U1277 (.IN1(n35), .IN2(n1545), .IN3(n1552), .IN4(n1), .Q(n1141));
   AO222X1 U1278 (.IN1(n464), .IN2(n1142), .IN3(n8), .IN4(n1143), .IN5(n1144), .IN6(n40), .
          Q(n1136));
   NAND3X0 U1279 (.IN1(n1145), .IN2(n420), .IN3(n1146), .QN(n1144));
   OA222X1 U1280 (.IN1(n1566), .IN2(n416), .IN3(n1568), .IN4(n332), .IN5(sboxw[1]), .IN6(
          n1542), .Q(n1146));
   OA22X1 U1281 (.IN1(n1567), .IN2(n1560), .IN3(n396), .IN4(n1555), .Q(n1145));
   NAND3X0 U1282 (.IN1(n442), .IN2(n478), .IN3(n352), .QN(n1143));
   AO221X1 U1283 (.IN1(n391), .IN2(n1569), .IN3(n15), .IN4(n411), .IN5(n1147), .Q(n1142)
          );
   AO22X1 U1284 (.IN1(n349), .IN2(n1568), .IN3(n447), .IN4(n1571), .Q(n1147));
   OA222X1 U1285 (.IN1(n1568), .IN2(n1549), .IN3(n1150), .IN4(n1571), .IN5(n7), .IN6(n679)
          , .Q(n1149));
   OA222X1 U1286 (.IN1(n1561), .IN2(n1), .IN3(n15), .IN4(n1558), .IN5(n331), .IN6(n1545), .
          Q(n1148));
   AO222X1 U1287 (.IN1(n917), .IN2(n1151), .IN3(n919), .IN4(n1152), .IN5(n1153), .IN6(n91)
          , .Q(new_sboxw[19]));
   AO221X1 U1288 (.IN1(n924), .IN2(n1154), .IN3(n922), .IN4(n1155), .IN5(n1156), .Q(n1153)
          );
   NAND3X0 U1290 (.IN1(n1159), .IN2(n1069), .IN3(n1160), .QN(n1158));
   OA22X1 U1291 (.IN1(n133), .IN2(n117), .IN3(n113), .IN4(n131), .Q(n1160));
   NAND3X0 U1292 (.IN1(n985), .IN2(n115), .IN3(n125), .QN(n1159));
   NAND4X0 U1293 (.IN1(n1161), .IN2(n1038), .IN3(n1162), .IN4(n1163), .QN(n1157));
   AOI222X1 U1294 (.IN1(n1062), .IN2(n1032), .IN3(n133), .IN4(n1048), .IN5(n1164), .IN6(
          n946), .QN(n1163));
   OA22X1 U1295 (.IN1(n128), .IN2(n44), .IN3(n132), .IN4(n22), .Q(n1032));
   OA22X1 U1296 (.IN1(n133), .IN2(n118), .IN3(n32), .IN4(n122), .Q(n1162));
   NAND4X0 U1297 (.IN1(n1096), .IN2(n114), .IN3(n1037), .IN4(n1165), .QN(n1155));
   OA222X1 U1298 (.IN1(n125), .IN2(n132), .IN3(n21), .IN4(n1095), .IN5(n985), .IN6(n118), .
          Q(n1165));
   NAND3X0 U1299 (.IN1(n23), .IN2(n128), .IN3(n31), .QN(n1096));
   NAND4X0 U1300 (.IN1(n967), .IN2(n1106), .IN3(n1167), .IN4(n1168), .QN(n1154));
   OA222X1 U1301 (.IN1(n1003), .IN2(n114), .IN3(n133), .IN4(n122), .IN5(n129), .IN6(n107)
          , .Q(n1168));
   NAND3X0 U1302 (.IN1(n131), .IN2(n115), .IN3(n125), .QN(n1167));
   NAND4X0 U1303 (.IN1(n1169), .IN2(n1170), .IN3(n1171), .IN4(n1172), .QN(n1152));
   OA222X1 U1304 (.IN1(n1173), .IN2(n45), .IN3(n10), .IN4(n1174), .IN5(n129), .IN6(n101), .
          Q(n1172));
   NOR4X0 U1305 (.IN1(n1175), .IN2(n1176), .IN3(n1177), .IN4(n1178), .QN(n1173));
   AO222X1 U1306 (.IN1(n1164), .IN2(n131), .IN3(n1048), .IN4(n31), .IN5(n1003), .IN6(n1062)
          , .Q(n1175));
   OA22X1 U1307 (.IN1(n21), .IN2(n22), .IN3(n132), .IN4(n128), .Q(n1003));
   NAND3X0 U1308 (.IN1(sboxw[17]), .IN2(n110), .IN3(n981), .QN(n1171));
   NAND3X0 U1309 (.IN1(n21), .IN2(n23), .IN3(n942), .QN(n1169));
   NAND4X0 U1310 (.IN1(n1170), .IN2(n1069), .IN3(n1179), .IN4(n1180), .QN(n1151));
   OA222X1 U1311 (.IN1(n1181), .IN2(n45), .IN3(n123), .IN4(n940), .IN5(n44), .IN6(n101), .
          Q(n1180));
   NOR4X0 U1312 (.IN1(n1182), .IN2(n1183), .IN3(n1184), .IN4(n1185), .QN(n1181));
   AO222X1 U1313 (.IN1(n1187), .IN2(n957), .IN3(n931), .IN4(n131), .IN5(n1001), .IN6(n130)
          , .Q(n1182));
   NAND3X0 U1314 (.IN1(n1025), .IN2(n45), .IN3(n1006), .QN(n1170));
   AO222X1 U1315 (.IN1(n917), .IN2(n1189), .IN3(n919), .IN4(n1190), .IN5(n1191), .IN6(n91)
          , .Q(new_sboxw[18]));
   AO221X1 U1316 (.IN1(n990), .IN2(n1192), .IN3(n924), .IN4(n1193), .IN5(n1194), .Q(n1191)
          );
   NAND4X0 U1318 (.IN1(n1007), .IN2(n1024), .IN3(n1197), .IN4(n1198), .QN(n1196));
   OA222X1 U1319 (.IN1(n1011), .IN2(n119), .IN3(sboxw[17]), .IN4(n108), .IN5(n31), .IN6(
          n122), .Q(n1198));
   OA22X1 U1320 (.IN1(n129), .IN2(n1114), .IN3(n128), .IN4(n1031), .Q(n1197));
   NAND4X0 U1321 (.IN1(n1024), .IN2(n1106), .IN3(n948), .IN4(n1199), .QN(n1195));
   OA22X1 U1322 (.IN1(n130), .IN2(n1200), .IN3(n132), .IN4(n1114), .Q(n1199));
   OA221X1 U1323 (.IN1(sboxw[17]), .IN2(n111), .IN3(n1203), .IN4(n132), .IN5(n1204), .Q(
          n1202));
   OA222X1 U1324 (.IN1(n109), .IN2(n32), .IN3(n957), .IN4(n122), .IN5(n129), .IN6(n120), .
          Q(n1201));
   NAND4X0 U1325 (.IN1(n1106), .IN2(n1093), .IN3(n1205), .IN4(n1206), .QN(n1192));
   OA221X1 U1326 (.IN1(n13), .IN2(n113), .IN3(n129), .IN4(n118), .IN5(n1207), .Q(n1206));
   AO221X1 U1327 (.IN1(n1208), .IN2(n44), .IN3(n10), .IN4(n1209), .IN5(n1210), .Q(n1190)
          );
   NAND3X0 U1328 (.IN1(n103), .IN2(n1211), .IN3(n1212), .QN(n1210));
   NAND3X0 U1329 (.IN1(n130), .IN2(n109), .IN3(n981), .QN(n1212));
   NAND4X0 U1330 (.IN1(n1213), .IN2(n121), .IN3(n1214), .IN4(n1215), .QN(n1209));
   NAND3X0 U1331 (.IN1(n956), .IN2(n32), .IN3(n23), .QN(n1213));
   AO221X1 U1332 (.IN1(n10), .IN2(n1216), .IN3(n1217), .IN4(n45), .IN5(n1218), .Q(n1189)
          );
   NAND4X0 U1334 (.IN1(n936), .IN2(n117), .IN3(n1219), .IN4(n1220), .QN(n1217));
   OA222X1 U1335 (.IN1(n129), .IN2(n111), .IN3(n1221), .IN4(n44), .IN5(n132), .IN6(n1095)
          , .Q(n1220));
   NAND3X0 U1336 (.IN1(n1222), .IN2(n1024), .IN3(n1207), .QN(n1216));
   OA22X1 U1337 (.IN1(n117), .IN2(n44), .IN3(n120), .IN4(n1011), .Q(n1207));
   AO22X1 U1338 (.IN1(sboxw[23]), .IN2(n1223), .IN3(n1224), .IN4(n91), .Q(new_sboxw[17])
          );
   AO222X1 U1339 (.IN1(n922), .IN2(n1225), .IN3(n924), .IN4(n1226), .IN5(n1227), .IN6(n92)
          , .Q(n1224));
   NAND4X0 U1340 (.IN1(n1228), .IN2(n941), .IN3(n1229), .IN4(n1230), .QN(n1227));
   OA221X1 U1341 (.IN1(n949), .IN2(n119), .IN3(n1116), .IN4(n100), .IN5(n1231), .Q(n1230)
          );
   OA22X1 U1342 (.IN1(n1011), .IN2(n94), .IN3(n130), .IN4(n101), .Q(n1231));
   OA22X1 U1343 (.IN1(n44), .IN2(n126), .IN3(n109), .IN4(n13), .Q(n1116));
   OA22X1 U1344 (.IN1(n128), .IN2(n31), .IN3(n985), .IN4(n22), .Q(n949));
   OA22X1 U1345 (.IN1(n1232), .IN2(n45), .IN3(n946), .IN4(n95), .Q(n1229));
   OA22X1 U1346 (.IN1(n133), .IN2(n107), .IN3(n31), .IN4(n113), .Q(n1232));
   NAND3X0 U1347 (.IN1(n133), .IN2(n45), .IN3(n1002), .QN(n1228));
   NAND4X0 U1348 (.IN1(n1092), .IN2(n951), .IN3(n1233), .IN4(n1234), .QN(n1226));
   OA222X1 U1349 (.IN1(n107), .IN2(n131), .IN3(n129), .IN4(n111), .IN5(n130), .IN6(n120), .
          Q(n1234));
   OA22X1 U1350 (.IN1(n946), .IN2(n1203), .IN3(n133), .IN4(n108), .Q(n1233));
   NAND4X0 U1351 (.IN1(n116), .IN2(n969), .IN3(n1235), .IN4(n1236), .QN(n1225));
   OA22X1 U1353 (.IN1(n133), .IN2(n1237), .IN3(n31), .IN4(n1090), .Q(n1235));
   AO221X1 U1354 (.IN1(n922), .IN2(n1238), .IN3(n1239), .IN4(n92), .IN5(n1240), .Q(n1223)
          );
   AO22X1 U1355 (.IN1(n924), .IN2(n1241), .IN3(n1242), .IN4(n932), .Q(n1240));
   NAND4X0 U1356 (.IN1(n1060), .IN2(n1091), .IN3(n1243), .IN4(n1244), .QN(n1241));
   OA22X1 U1357 (.IN1(n31), .IN2(n107), .IN3(n114), .IN4(n32), .Q(n1244));
   AO222X1 U1358 (.IN1(n1079), .IN2(n1245), .IN3(n10), .IN4(n1246), .IN5(n1247), .IN6(n45)
          , .Q(n1239));
   NAND3X0 U1359 (.IN1(n1248), .IN2(n1035), .IN3(n1249), .QN(n1247));
   OA222X1 U1360 (.IN1(n128), .IN2(n1031), .IN3(n130), .IN4(n947), .IN5(sboxw[17]), .IN6(
          n104), .Q(n1249));
   OA22X1 U1361 (.IN1(n129), .IN2(n122), .IN3(n1011), .IN4(n117), .Q(n1248));
   NAND3X0 U1362 (.IN1(n1057), .IN2(n1093), .IN3(n967), .QN(n1246));
   AO221X1 U1363 (.IN1(n1006), .IN2(n131), .IN3(n21), .IN4(n1026), .IN5(n1250), .Q(n1245)
          );
   AO22X1 U1364 (.IN1(n964), .IN2(n130), .IN3(n1062), .IN4(n133), .Q(n1250));
   OA222X1 U1365 (.IN1(n130), .IN2(n111), .IN3(n1253), .IN4(n133), .IN5(n957), .IN6(n1203)
          , .Q(n1252));
   OA222X1 U1366 (.IN1(n123), .IN2(n32), .IN3(n21), .IN4(n120), .IN5(n946), .IN6(n107), .Q(
          n1251));
   AO22X1 U1367 (.IN1(sboxw[23]), .IN2(n1254), .IN3(n1255), .IN4(n91), .Q(new_sboxw[16])
          );
   NAND4X0 U1369 (.IN1(n1258), .IN2(n98), .IN3(n1259), .IN4(n1260), .QN(n1257));
   AOI222X1 U1370 (.IN1(n10), .IN2(n1261), .IN3(n1262), .IN4(n45), .IN5(n1075), .IN6(n44)
          , .QN(n1260));
   NAND3X0 U1371 (.IN1(n961), .IN2(n968), .IN3(n1263), .QN(n1262));
   NAND4X0 U1372 (.IN1(n1057), .IN2(n117), .IN3(n1265), .IN4(n1266), .QN(n1261));
   OA222X1 U1373 (.IN1(n133), .IN2(n119), .IN3(n130), .IN4(n1095), .IN5(n32), .IN6(n111), .
          Q(n1266));
   OR2X1 U1374 (.IN1(n1114), .IN2(n133), .Q(n1204));
   NAND3X0 U1375 (.IN1(n31), .IN2(n23), .IN3(n942), .QN(n1258));
   NAND4X0 U1376 (.IN1(n1268), .IN2(n1211), .IN3(n1269), .IN4(n1270), .QN(n1256));
   AOI222X1 U1377 (.IN1(n10), .IN2(n1271), .IN3(n1055), .IN4(n131), .IN5(n1075), .IN6(n132)
          , .QN(n1270));
   NAND4X0 U1378 (.IN1(n1219), .IN2(n1093), .IN3(n1272), .IN4(n1273), .QN(n1271));
   OA222X1 U1379 (.IN1(n1011), .IN2(n113), .IN3(n31), .IN4(n118), .IN5(n985), .IN6(n120), .
          Q(n1273));
   NAND3X0 U1380 (.IN1(n131), .IN2(n128), .IN3(n110), .QN(n1219));
   AO222X1 U1382 (.IN1(sboxw[22]), .IN2(n1274), .IN3(n922), .IN4(n1275), .IN5(n1276), .IN6(
          n92), .Q(n1254));
   AO221X1 U1383 (.IN1(n1277), .IN2(n45), .IN3(n1001), .IN4(n985), .IN5(n1278), .Q(n1276)
          );
   AO222X1 U1384 (.IN1(n974), .IN2(n132), .IN3(n1279), .IN4(n22), .IN5(n981), .IN6(n1280)
          , .Q(n1278));
   AO221X1 U1385 (.IN1(n957), .IN2(n1062), .IN3(n1006), .IN4(n133), .IN5(n1061), .Q(n1280)
          );
   AO221X1 U1387 (.IN1(n985), .IN2(n1002), .IN3(n964), .IN4(n1264), .IN5(n971), .Q(n1275)
          );
   XNOR2X1 U1388 (.IN1(n22), .IN2(n21), .Q(n1282));
   AO221X1 U1389 (.IN1(n1283), .IN2(n1011), .IN3(n10), .IN4(n1284), .IN5(n1188), .Q(n1274)
          );
   NAND4X0 U1390 (.IN1(n112), .IN2(n111), .IN3(n1285), .IN4(n1286), .QN(n1284));
   OA221X1 U1391 (.IN1(n13), .IN2(n117), .IN3(n107), .IN4(n131), .IN5(n1287), .Q(n1286));
   OA22X1 U1392 (.IN1(n985), .IN2(n122), .IN3(n133), .IN4(n120), .Q(n1287));
   AO222X1 U1394 (.IN1(n188), .IN2(n1293), .IN3(n190), .IN4(n1294), .IN5(n1295), .IN6(n135)
          , .Q(n1292));
   NAND4X0 U1395 (.IN1(n1296), .IN2(n1297), .IN3(n1298), .IN4(n1299), .QN(n1295));
   NAND4X0 U1397 (.IN1(n1302), .IN2(n1303), .IN3(n1304), .IN4(n1305), .QN(n1301));
   OA22X1 U1398 (.IN1(n37), .IN2(n1306), .IN3(n148), .IN4(n1307), .Q(n1298));
   NAND3X0 U1399 (.IN1(n211), .IN2(n167), .IN3(n271), .QN(n1296));
   NAND4X0 U1400 (.IN1(n171), .IN2(n1308), .IN3(n1309), .IN4(n1310), .QN(n1294));
   OA222X1 U1401 (.IN1(n204), .IN2(n147), .IN3(n177), .IN4(n237), .IN5(n38), .IN6(n146), .
          Q(n1310));
   AND2X1 U1402 (.IN1(n157), .IN2(n1311), .Q(n1309));
   OA22X1 U1403 (.IN1(n281), .IN2(n19), .IN3(n172), .IN4(n38), .Q(n197));
   NAND4X0 U1404 (.IN1(n1312), .IN2(n207), .IN3(n1313), .IN4(n1314), .QN(n1293));
   OA22X1 U1405 (.IN1(n1315), .IN2(n177), .IN3(n176), .IN4(n157), .Q(n1314));
   NAND3X0 U1406 (.IN1(n1316), .IN2(n174), .IN3(n20), .QN(n1313));
   NAND3X0 U1407 (.IN1(n19), .IN2(n153), .IN3(n37), .QN(n1312));
   NAND4X0 U1408 (.IN1(n1317), .IN2(n1318), .IN3(n1319), .IN4(n1320), .QN(n1291));
   AOI222X1 U1409 (.IN1(n260), .IN2(n211), .IN3(n1321), .IN4(n43), .IN5(n9), .IN6(n1322), .
          QN(n1320));
   OAI221X1 U1410 (.IN1(n163), .IN2(n38), .IN3(n173), .IN4(n148), .IN5(n1308), .QN(n1322)
          );
   NAND3X0 U1411 (.IN1(n213), .IN2(n151), .IN3(n240), .QN(n1321));
   OA22X1 U1412 (.IN1(n41), .IN2(n137), .IN3(n1323), .IN4(n143), .Q(n1319));
   AND3X1 U1413 (.IN1(n1303), .IN2(n1324), .IN3(n1325), .Q(n1323));
   NAND3X0 U1414 (.IN1(n204), .IN2(n167), .IN3(n229), .QN(n1317));
   OA221X1 U1415 (.IN1(n147), .IN2(n1307), .IN3(n20), .IN4(n1328), .IN5(n1329), .Q(n1327)
          );
   OA22X1 U1416 (.IN1(n204), .IN2(n140), .IN3(n175), .IN4(n143), .Q(n1328));
   OA222X1 U1417 (.IN1(n1330), .IN2(n43), .IN3(n9), .IN4(n1331), .IN5(n143), .IN6(n1325), .
          Q(n1326));
   AND3X1 U1418 (.IN1(n1332), .IN2(n1333), .IN3(n1334), .Q(n1330));
   OA222X1 U1419 (.IN1(n161), .IN2(n281), .IN3(n237), .IN4(n38), .IN5(n176), .IN6(n146), .
          Q(n1332));
   AO22X1 U1420 (.IN1(n1335), .IN2(n134), .IN3(sboxw[15]), .IN4(n1336), .Q(new_sboxw[14])
          );
   AO222X1 U1421 (.IN1(n1337), .IN2(n1338), .IN3(n1339), .IN4(n1340), .IN5(sboxw[14]), .
          IN6(n1341), .Q(n1336));
   AO221X1 U1422 (.IN1(n9), .IN2(n1342), .IN3(n1343), .IN4(n43), .IN5(n1344), .Q(n1341));
   AO22X1 U1423 (.IN1(n223), .IN2(n38), .IN3(n200), .IN4(n204), .Q(n1344));
   OA222X1 U1424 (.IN1(n150), .IN2(n174), .IN3(n18), .IN4(n1347), .IN5(n165), .IN6(n176), .
          Q(n1346));
   OA222X1 U1425 (.IN1(n1350), .IN2(n148), .IN3(n158), .IN4(n3), .IN5(n163), .IN6(n175), .
          Q(n1345));
   NAND3X0 U1426 (.IN1(n1351), .IN2(n151), .IN3(n1352), .QN(n1342));
   AO221X1 U1428 (.IN1(n1354), .IN2(n177), .IN3(n1355), .IN4(n173), .IN5(n301), .Q(n1353)
          );
   NAND4X0 U1429 (.IN1(n1311), .IN2(n146), .IN3(n1356), .IN4(n1357), .QN(n1338));
   OA222X1 U1430 (.IN1(n41), .IN2(n148), .IN3(n211), .IN4(n152), .IN5(n158), .IN6(n174), .
          Q(n1357));
   OA22X1 U1431 (.IN1(n245), .IN2(n267), .IN3(n175), .IN4(n157), .Q(n1356));
   AO221X1 U1432 (.IN1(n188), .IN2(n1358), .IN3(n1359), .IN4(n135), .IN5(n1360), .Q(n1335)
          );
   AO22X1 U1433 (.IN1(n270), .IN2(sboxw[14]), .IN3(n190), .IN4(n1361), .Q(n1360));
   NAND3X0 U1434 (.IN1(n297), .IN2(n1362), .IN3(n1363), .QN(n1361));
   OA221X1 U1435 (.IN1(n18), .IN2(n150), .IN3(n3), .IN4(n145), .IN5(n1364), .Q(n1363));
   OA22X1 U1436 (.IN1(n173), .IN2(n148), .IN3(n158), .IN4(n41), .Q(n297));
   OA221X1 U1437 (.IN1(n1369), .IN2(n138), .IN3(n1370), .IN4(n140), .IN5(n1371), .Q(n1368)
          );
   AND2X1 U1438 (.IN1(n1303), .IN2(n236), .Q(n1369));
   OA222X1 U1439 (.IN1(n1372), .IN2(n159), .IN3(n1373), .IN4(n43), .IN5(n9), .IN6(n1374), .
          Q(n1367));
   OA22X1 U1440 (.IN1(n1372), .IN2(n148), .IN3(sboxw[11]), .IN4(n281), .Q(n1374));
   NAND4X0 U1441 (.IN1(n234), .IN2(n1376), .IN3(n1377), .IN4(n282), .QN(n1358));
   OR2X1 U1442 (.IN1(n163), .IN2(n1350), .Q(n1376));
   AO222X1 U1443 (.IN1(n1290), .IN2(n1378), .IN3(n1379), .IN4(n134), .IN5(n1288), .IN6(
          n1380), .Q(new_sboxw[13]));
   AO222X1 U1444 (.IN1(n286), .IN2(n1381), .IN3(n1382), .IN4(n43), .IN5(n9), .IN6(n1383), .
          Q(n1380));
   NAND4X0 U1445 (.IN1(n1308), .IN2(n1305), .IN3(n1384), .IN4(n1385), .QN(n1383));
   OA222X1 U1446 (.IN1(n159), .IN2(n175), .IN3(n1386), .IN4(n173), .IN5(n161), .IN6(n3), .
          Q(n1385));
   NAND3X0 U1447 (.IN1(n1331), .IN2(n1304), .IN3(n1387), .QN(n1382));
   AO221X1 U1448 (.IN1(n20), .IN2(n173), .IN3(n155), .IN4(n177), .IN5(n167), .Q(n1381));
   AO22X1 U1449 (.IN1(n1388), .IN2(n135), .IN3(sboxw[14]), .IN4(n1389), .Q(n1379));
   AO221X1 U1450 (.IN1(n286), .IN2(n1390), .IN3(n9), .IN4(n1391), .IN5(n1392), .Q(n1389)
          );
   AO22X1 U1451 (.IN1(n277), .IN2(n18), .IN3(n1393), .IN4(n271), .Q(n1392));
   NAND4X0 U1452 (.IN1(n1384), .IN2(n160), .IN3(n1394), .IN4(n1395), .QN(n1391));
   OA221X1 U1453 (.IN1(n29), .IN2(n146), .IN3(n42), .IN4(n157), .IN5(n224), .Q(n1395));
   AND2X1 U1454 (.IN1(n238), .IN2(n151), .Q(n1394));
   OR2X1 U1455 (.IN1(n237), .IN2(n176), .Q(n1384));
   AO222X1 U1456 (.IN1(n30), .IN2(n245), .IN3(n37), .IN4(n241), .IN5(n244), .IN6(n176), .Q(
          n1390));
   NAND4X0 U1457 (.IN1(n214), .IN2(n238), .IN3(n1396), .IN4(n1397), .QN(n1388));
   OA221X1 U1458 (.IN1(n1398), .IN2(n43), .IN3(n9), .IN4(n1399), .IN5(n1400), .Q(n1397));
   OA22X1 U1459 (.IN1(n1401), .IN2(n138), .IN3(n28), .IN4(n157), .Q(n1400));
   AND3X1 U1460 (.IN1(n236), .IN2(n163), .IN3(n1331), .Q(n1401));
   NAND4X0 U1461 (.IN1(n1297), .IN2(n207), .IN3(n1404), .IN4(n1405), .QN(n1378));
   OA222X1 U1462 (.IN1(n1406), .IN2(n43), .IN3(n9), .IN4(n1407), .IN5(n3), .IN6(n142), .Q(
          n1405));
   OA22X1 U1463 (.IN1(n152), .IN2(n41), .IN3(n174), .IN4(n162), .Q(n1334));
   OA221X1 U1464 (.IN1(n163), .IN2(n42), .IN3(n38), .IN4(n147), .IN5(n1408), .Q(n1406));
   OA22X1 U1465 (.IN1(n138), .IN2(n1409), .IN3(n1410), .IN4(n143), .Q(n1404));
   NAND3X0 U1466 (.IN1(n245), .IN2(n3), .IN3(n229), .QN(n1297));
   AO22X1 U1467 (.IN1(n1411), .IN2(n134), .IN3(sboxw[15]), .IN4(n1412), .Q(new_sboxw[12])
          );
   AO222X1 U1468 (.IN1(n1337), .IN2(n1413), .IN3(n1339), .IN4(n1414), .IN5(sboxw[14]), .
          IN6(n1415), .Q(n1412));
   OAI222X1 U1469 (.IN1(n1416), .IN2(n43), .IN3(n1417), .IN4(n138), .IN5(n9), .IN6(n1418)
          , .QN(n1415));
   OAI222X1 U1470 (.IN1(n150), .IN2(n38), .IN3(n217), .IN4(n204), .IN5(n157), .IN6(n41), .
          QN(n1420));
   NAND4X0 U1471 (.IN1(n225), .IN2(n1304), .IN3(n208), .IN4(n239), .QN(n1419));
   OA221X1 U1472 (.IN1(n148), .IN2(n176), .IN3(n175), .IN4(n145), .IN5(n1421), .Q(n1416)
          );
   NAND4X0 U1473 (.IN1(n1422), .IN2(n239), .IN3(n1423), .IN4(n1424), .QN(n1414));
   OA222X1 U1474 (.IN1(n204), .IN2(n162), .IN3(n42), .IN4(n217), .IN5(n173), .IN6(n157), .
          Q(n1424));
   NAND3X0 U1475 (.IN1(n19), .IN2(n173), .IN3(n266), .QN(n1423));
   NAND3X0 U1476 (.IN1(n1352), .IN2(n1425), .IN3(n1426), .QN(n1413));
   OA221X1 U1477 (.IN1(n161), .IN2(n176), .IN3(n150), .IN4(n173), .IN5(n1427), .Q(n1426)
          );
   NAND3X0 U1478 (.IN1(n174), .IN2(n172), .IN3(n266), .QN(n1427));
   OA22X1 U1479 (.IN1(n162), .IN2(n30), .IN3(n145), .IN4(n176), .Q(n1352));
   AO221X1 U1480 (.IN1(n1337), .IN2(n1428), .IN3(sboxw[14]), .IN4(n1429), .IN5(n1430), .Q(
          n1411));
   AO22X1 U1481 (.IN1(n1339), .IN2(n1431), .IN3(n281), .IN4(n200), .Q(n1430));
   NAND4X0 U1482 (.IN1(n1432), .IN2(n1305), .IN3(n1433), .IN4(n1434), .QN(n1431));
   OA222X1 U1483 (.IN1(n146), .IN2(n176), .IN3(n175), .IN4(n164), .IN5(n204), .IN6(n157), .
          Q(n1434));
   NAND3X0 U1484 (.IN1(n154), .IN2(n173), .IN3(n19), .QN(n1433));
   AO222X1 U1485 (.IN1(n1435), .IN2(n43), .IN3(n286), .IN4(n1436), .IN5(n9), .IN6(n1437), .
          Q(n1429));
   NAND4X0 U1486 (.IN1(n156), .IN2(n145), .IN3(n1438), .IN4(n1439), .QN(n1437));
   OA222X1 U1487 (.IN1(n153), .IN2(n175), .IN3(n173), .IN4(n169), .IN5(n161), .IN6(n177), .
          Q(n1439));
   AO21X1 U1488 (.IN1(n148), .IN2(n166), .IN3(n37), .Q(n1438));
   NAND3X0 U1489 (.IN1(n1441), .IN2(n163), .IN3(n198), .QN(n1436));
   OA22X1 U1490 (.IN1(n42), .IN2(n167), .IN3(n153), .IN4(n41), .Q(n198));
   OAI221X1 U1491 (.IN1(n152), .IN2(n204), .IN3(n147), .IN4(n173), .IN5(n208), .QN(n1435)
          );
   NAND4X0 U1492 (.IN1(n1308), .IN2(n162), .IN3(n1442), .IN4(n1443), .QN(n1428));
   OA22X1 U1493 (.IN1(n163), .IN2(n174), .IN3(n38), .IN4(n159), .Q(n1443));
   AO222X1 U1494 (.IN1(n1288), .IN2(n1444), .IN3(n1290), .IN4(n1445), .IN5(n1446), .IN6(
          n134), .Q(new_sboxw[11]));
   AO221X1 U1495 (.IN1(n1337), .IN2(n1447), .IN3(n1339), .IN4(n1448), .IN5(n1449), .Q(
          n1446));
   AO22X1 U1496 (.IN1(n188), .IN2(n1450), .IN3(n190), .IN4(n1451), .Q(n1449));
   NAND4X0 U1497 (.IN1(n1452), .IN2(n1432), .IN3(n1453), .IN4(n1454), .QN(n1451));
   OA222X1 U1498 (.IN1(n211), .IN2(n152), .IN3(n161), .IN4(n177), .IN5(n18), .IN6(n146), .
          Q(n1454));
   NAND3X0 U1499 (.IN1(n175), .IN2(n155), .IN3(n168), .QN(n1452));
   NAND4X0 U1500 (.IN1(n1422), .IN2(n148), .IN3(n1377), .IN4(n1455), .QN(n1450));
   OA222X1 U1501 (.IN1(n159), .IN2(n170), .IN3(n18), .IN4(n265), .IN5(n217), .IN6(n176), .
          Q(n1455));
   NAND4X0 U1502 (.IN1(n1456), .IN2(n282), .IN3(n1457), .IN4(n1458), .QN(n1448));
   OA222X1 U1503 (.IN1(n153), .IN2(n170), .IN3(n18), .IN4(n162), .IN5(n175), .IN6(n147), .
          Q(n1458));
   OA22X1 U1504 (.IN1(n42), .IN2(n172), .IN3(n176), .IN4(n19), .Q(n1372));
   OA22X1 U1505 (.IN1(n177), .IN2(n157), .IN3(n146), .IN4(n174), .Q(n1457));
   NAND3X0 U1506 (.IN1(n1459), .IN2(n1402), .IN3(n1460), .QN(n1447));
   OA22X1 U1507 (.IN1(n158), .IN2(n177), .IN3(n175), .IN4(n147), .Q(n1460));
   NAND3X0 U1508 (.IN1(n281), .IN2(n155), .IN3(n168), .QN(n1459));
   NAND4X0 U1509 (.IN1(n1461), .IN2(n1462), .IN3(n1463), .IN4(n1464), .QN(n1445));
   OA222X1 U1510 (.IN1(n1465), .IN2(n43), .IN3(n9), .IN4(n1466), .IN5(n211), .IN6(n139), .
          Q(n1464));
   AO222X1 U1511 (.IN1(n1375), .IN2(n175), .IN3(n37), .IN4(n228), .IN5(n1350), .IN6(n241)
          , .Q(n1468));
   OA22X1 U1512 (.IN1(n19), .IN2(n18), .IN3(n176), .IN4(n172), .Q(n1350));
   AO222X1 U1513 (.IN1(n1348), .IN2(n28), .IN3(n211), .IN4(n1469), .IN5(n1470), .IN6(n41)
          , .Q(n1467));
   NAND3X0 U1515 (.IN1(n18), .IN2(n20), .IN3(n271), .QN(n1461));
   NAND4X0 U1516 (.IN1(n1462), .IN2(n1402), .IN3(n1471), .IN4(n1472), .QN(n1444));
   OA222X1 U1517 (.IN1(n1473), .IN2(n43), .IN3(n163), .IN4(n1307), .IN5(n42), .IN6(n139), .
          Q(n1472));
   AO222X1 U1518 (.IN1(n1300), .IN2(n175), .IN3(n1470), .IN4(n174), .IN5(n1375), .IN6(n30)
          , .Q(n1475));
   NAND3X0 U1520 (.IN1(n1365), .IN2(n43), .IN3(n245), .QN(n1462));
   AO221X1 U1522 (.IN1(n1339), .IN2(n1479), .IN3(n190), .IN4(n1480), .IN5(n1481), .Q(n1478)
          );
   AO22X1 U1523 (.IN1(n188), .IN2(n1482), .IN3(n1337), .IN4(n1483), .Q(n1481));
   NAND4X0 U1524 (.IN1(n1484), .IN2(n1364), .IN3(n1485), .IN4(n1486), .QN(n1483));
   OA222X1 U1525 (.IN1(n28), .IN2(n159), .IN3(n41), .IN4(n150), .IN5(n38), .IN6(n161), .Q(
          n1486));
   OA22X1 U1526 (.IN1(n211), .IN2(n169), .IN3(n172), .IN4(n236), .Q(n1485));
   NAND4X0 U1527 (.IN1(n1364), .IN2(n1432), .IN3(n1311), .IN4(n1487), .QN(n1482));
   OA22X1 U1528 (.IN1(n173), .IN2(n1488), .IN3(n176), .IN4(n169), .Q(n1487));
   OA221X1 U1529 (.IN1(n161), .IN2(n174), .IN3(n212), .IN4(n176), .IN5(n268), .Q(n1490));
   OA222X1 U1530 (.IN1(n153), .IN2(n3), .IN3(n41), .IN4(n146), .IN5(n211), .IN6(n162), .Q(
          n1489));
   NAND4X0 U1531 (.IN1(n1432), .IN2(n239), .IN3(n1491), .IN4(n1492), .QN(n1479));
   OA221X1 U1532 (.IN1(n41), .IN2(n147), .IN3(n28), .IN4(n146), .IN5(n1493), .Q(n1492));
   AO221X1 U1533 (.IN1(n202), .IN2(n42), .IN3(n9), .IN4(n1494), .IN5(n1495), .Q(n1477));
   NAND3X0 U1534 (.IN1(n141), .IN2(n273), .IN3(n1496), .QN(n1495));
   NAND3X0 U1535 (.IN1(n153), .IN2(n173), .IN3(n286), .QN(n1496));
   NAND4X0 U1537 (.IN1(n1497), .IN2(n1371), .IN3(n1498), .IN4(n1499), .QN(n1494));
   NAND3X0 U1538 (.IN1(n1316), .IN2(n3), .IN3(n20), .QN(n1497));
   AO221X1 U1539 (.IN1(n9), .IN2(n1500), .IN3(n1501), .IN4(n43), .IN5(n1502), .Q(n1476));
   AO221X1 U1540 (.IN1(n290), .IN2(n211), .IN3(n223), .IN4(n174), .IN5(n136), .Q(n1502));
   NAND4X0 U1541 (.IN1(n1305), .IN2(n158), .IN3(n278), .IN4(n1503), .QN(n1501));
   NAND3X0 U1543 (.IN1(n175), .IN2(n172), .IN3(n154), .QN(n278));
   NAND3X0 U1544 (.IN1(n1505), .IN2(n1364), .IN3(n1493), .QN(n1500));
   OA22X1 U1545 (.IN1(n42), .IN2(n158), .IN3(n162), .IN4(n29), .Q(n1493));
   AO22X1 U1547 (.IN1(n1508), .IN2(n179), .IN3(sboxw[6]), .IN4(n1509), .Q(n1507));
   NAND4X0 U1548 (.IN1(n1510), .IN2(n185), .IN3(n1511), .IN4(n1512), .QN(n1509));
   NAND3X0 U1550 (.IN1(n346), .IN2(n353), .IN3(n1515), .QN(n1514));
   NAND4X0 U1551 (.IN1(n442), .IN2(n1555), .IN3(n1517), .IN4(n1518), .QN(n1513));
   OA222X1 U1552 (.IN1(n1571), .IN2(n1557), .IN3(n1568), .IN4(n480), .IN5(n1), .IN6(n1549)
          , .Q(n1518));
   OR2X1 U1553 (.IN1(n499), .IN2(n1571), .Q(n680));
   NAND3X0 U1554 (.IN1(n35), .IN2(n17), .IN3(n327), .QN(n1510));
   NAND4X0 U1555 (.IN1(n1520), .IN2(n687), .IN3(n1521), .IN4(n1522), .QN(n1508));
   NAND4X0 U1557 (.IN1(n695), .IN2(n478), .IN3(n1524), .IN4(n1525), .QN(n1523));
   OA222X1 U1558 (.IN1(n396), .IN2(n1551), .IN3(n36), .IN4(n1556), .IN5(n370), .IN6(n1558)
          , .Q(n1525));
   NAND3X0 U1559 (.IN1(n1569), .IN2(n1566), .IN3(n1548), .QN(n695));
   NAND3X0 U1560 (.IN1(n7), .IN2(n1548), .IN3(n327), .QN(n1520));
   AO222X1 U1561 (.IN1(sboxw[6]), .IN2(n1526), .IN3(n307), .IN4(n1527), .IN5(n1528), .IN6(
          n179), .Q(n1506));
   AO221X1 U1562 (.IN1(n1529), .IN2(n40), .IN3(n386), .IN4(n370), .IN5(n1530), .Q(n1528)
          );
   AO222X1 U1563 (.IN1(n359), .IN2(n1570), .IN3(n1531), .IN4(n16), .IN5(n366), .IN6(n1532)
          , .Q(n1530));
   AO221X1 U1564 (.IN1(n342), .IN2(n447), .IN3(n391), .IN4(n1571), .IN5(n446), .Q(n1532)
          );
   OAI221X1 U1565 (.IN1(n1558), .IN2(n331), .IN3(n1555), .IN4(n396), .IN5(n476), .QN(n1529)
          );
   AO221X1 U1566 (.IN1(n370), .IN2(n387), .IN3(n349), .IN4(n1516), .IN5(n356), .Q(n1527)
          );
   XNOR2X1 U1567 (.IN1(n16), .IN2(n15), .Q(n1534));
   AO221X1 U1568 (.IN1(n1535), .IN2(n396), .IN3(n8), .IN4(n1536), .IN5(n542), .Q(n1526));
   NAND4X0 U1569 (.IN1(n1550), .IN2(n1549), .IN3(n1537), .IN4(n1538), .QN(n1536));
   OA221X1 U1570 (.IN1(n12), .IN2(n1555), .IN3(n1545), .IN4(n1569), .IN5(n1539), .Q(n1538)
          );
   OA22X1 U1571 (.IN1(n370), .IN2(n1560), .IN3(n1571), .IN4(n1558), .Q(n1539));
   NBUFFX2 U1 (.INP(sboxw[16]), .Z(n21));
   NBUFFX2 U2 (.INP(sboxw[18]), .Z(n22));
   NBUFFX2 U3 (.INP(sboxw[8]), .Z(n18));
   NBUFFX2 U4 (.INP(sboxw[24]), .Z(n24));
   NBUFFX2 U5 (.INP(sboxw[12]), .Z(n20));
   NBUFFX2 U6 (.INP(sboxw[26]), .Z(n25));
   NBUFFX2 U7 (.INP(sboxw[2]), .Z(n16));
   NBUFFX2 U8 (.INP(sboxw[0]), .Z(n15));
   NBUFFX2 U9 (.INP(sboxw[10]), .Z(n19));
   INVX0 U10 (.INP(n1185), .ZN(n116));
   INVX0 U11 (.INP(n539), .ZN(n1554));
   OA21X1 U12 (.IN1(n89), .IN2(n56), .IN3(n604), .Q(n808));
   INVX0 U13 (.INP(n814), .ZN(n73));
   OA21X1 U14 (.IN1(n132), .IN2(n99), .IN3(n978), .Q(n1179));
   NOR2X0 U15 (.IN1(n1061), .IN2(n1047), .QN(n1058));
   INVX0 U16 (.INP(n370), .ZN(n1570));
   NOR2X0 U17 (.IN1(n446), .IN2(n432), .QN(n443));
   INVX0 U18 (.INP(n611), .ZN(n89));
   NOR2X0 U19 (.IN1(n721), .IN2(n707), .QN(n718));
   NOR2X0 U20 (.IN1(n117), .IN2(n31), .QN(n1185));
   INVX0 U21 (.INP(n972), .ZN(n105));
   NOR2X0 U22 (.IN1(n1555), .IN2(n35), .QN(n539));
   INVX0 U23 (.INP(n538), .ZN(n1550));
   INVX0 U24 (.INP(n980), .ZN(n106));
   INVX0 U25 (.INP(n301), .ZN(n156));
   INVX0 U26 (.INP(n1177), .ZN(n121));
   INVX0 U27 (.INP(n1184), .ZN(n112));
   INVX0 U28 (.INP(n813), .ZN(n69));
   NOR2X0 U29 (.IN1(n74), .IN2(n33), .QN(n814));
   INVX0 U30 (.INP(n806), .ZN(n78));
   INVX0 U31 (.INP(n531), .ZN(n1559));
   INVX0 U32 (.INP(n622), .ZN(n51));
   INVX0 U33 (.INP(n365), .ZN(n1544));
   INVX0 U34 (.INP(n357), .ZN(n1543));
   INVX0 U35 (.INP(n606), .ZN(n63));
   NAND2X1 U36 (.IN1(n817), .IN2(n33), .QN(n604));
   INVX0 U37 (.INP(n598), .ZN(n62));
   NAND2X1 U38 (.IN1(n1188), .IN2(n938), .QN(n978));
   INVX0 U39 (.INP(n896), .ZN(n56));
   INVX0 U40 (.INP(n1267), .ZN(n99));
   INVX0 U41 (.INP(n290), .ZN(n137));
   INVX0 U42 (.INP(n974), .ZN(n95));
   INVX0 U43 (.INP(n1075), .ZN(n97));
   INVX0 U44 (.INP(n260), .ZN(n142));
   INVX0 U45 (.INP(n735), .ZN(n54));
   INVX0 U46 (.INP(n270), .ZN(n144));
   INVX0 U47 (.INP(n1), .ZN(n35));
   INVX0 U48 (.INP(n342), .ZN(n1567));
   NAND2X1 U49 (.IN1(n433), .IN2(n1567), .QN(n1140));
   NOR2X0 U50 (.IN1(n1571), .IN2(n12), .QN(n370));
   NOR2X0 U51 (.IN1(n332), .IN2(n1570), .QN(n432));
   OA21X1 U52 (.IN1(sboxw[1]), .IN2(n1558), .IN3(n354), .Q(n418));
   NOR2X0 U53 (.IN1(n90), .IN2(n14), .QN(n611));
   NOR2X0 U54 (.IN1(n573), .IN2(n89), .QN(n707));
   NAND2X1 U55 (.IN1(n1569), .IN2(n401), .QN(n410));
   OA21X1 U56 (.IN1(n985), .IN2(n123), .IN3(n1069), .Q(n1066));
   OA21X1 U57 (.IN1(n370), .IN2(n1561), .IN3(n454), .Q(n451));
   INVX0 U58 (.INP(n938), .ZN(n32));
   NAND2X1 U59 (.IN1(n387), .IN2(n1569), .QN(n502));
   NOR2X0 U60 (.IN1(n31), .IN2(n955), .QN(n1056));
   NAND2X1 U61 (.IN1(n88), .IN2(n642), .QN(n651));
   NAND2X1 U62 (.IN1(n1201), .IN2(n1202), .QN(n1193));
   NAND2X1 U63 (.IN1(n1048), .IN2(n985), .QN(n935));
   NAND2X1 U64 (.IN1(n677), .IN2(n678), .QN(n669));
   INVX0 U65 (.INP(n583), .ZN(n86));
   NAND2X1 U66 (.IN1(n708), .IN2(n86), .QN(n872));
   NAND2X1 U67 (.IN1(n322), .IN2(n6), .QN(n423));
   AO221X1 U68 (.IN1(n974), .IN2(n129), .IN3(n932), .IN4(n957), .IN5(n973), .Q(n1218));
   NOR2X0 U69 (.IN1(n133), .IN2(n109), .QN(n972));
   NAND2X1 U70 (.IN1(n518), .IN2(n7), .QN(n442));
   OA21X1 U71 (.IN1(sboxw[25]), .IN2(n77), .IN3(n595), .Q(n659));
   NAND2X1 U72 (.IN1(n985), .IN2(n937), .QN(n967));
   OA21X1 U73 (.IN1(n611), .IN2(n80), .IN3(n729), .Q(n726));
   INVX0 U74 (.INP(n411), .ZN(n1552));
   INVX0 U75 (.INP(n518), .ZN(n1551));
   NOR2X0 U76 (.IN1(n1568), .IN2(n1551), .QN(n538));
   NOR2X0 U77 (.IN1(n130), .IN2(n109), .QN(n980));
   NAND2X1 U78 (.IN1(n628), .IN2(n88), .QN(n777));
   NOR2X0 U79 (.IN1(n123), .IN2(n133), .QN(n1061));
   NOR2X0 U80 (.IN1(n281), .IN2(n27), .QN(n211));
   NOR2X0 U81 (.IN1(n157), .IN2(n174), .QN(n301));
   NAND2X1 U82 (.IN1(n1375), .IN2(n211), .QN(n213));
   NAND2X1 U83 (.IN1(n250), .IN2(n174), .QN(n282));
   OA21X1 U84 (.IN1(n37), .IN2(n157), .IN3(n282), .Q(n279));
   INVX0 U85 (.INP(n244), .ZN(n148));
   NAND2X1 U86 (.IN1(n937), .IN2(n133), .QN(n1092));
   NAND2X1 U87 (.IN1(n211), .IN2(n206), .QN(n1402));
   OA21X1 U88 (.IN1(n281), .IN2(n163), .IN3(n1402), .Q(n1399));
   NAND2X1 U89 (.IN1(n433), .IN2(n370), .QN(n320));
   NOR2X0 U90 (.IN1(n35), .IN2(n340), .QN(n441));
   INVX0 U91 (.INP(n2), .ZN(n33));
   NAND2X1 U92 (.IN1(n1375), .IN2(n174), .QN(n238));
   NAND2X1 U93 (.IN1(n1164), .IN2(n133), .QN(n936));
   NOR2X0 U94 (.IN1(n122), .IN2(n130), .QN(n1177));
   INVX0 U95 (.INP(n206), .ZN(n152));
   NAND2X1 U96 (.IN1(n830), .IN2(n831), .QN(n822));
   NOR2X0 U97 (.IN1(n130), .IN2(n113), .QN(n1184));
   INVX0 U98 (.INP(n1026), .ZN(n114));
   NAND2X1 U99 (.IN1(n708), .IN2(n611), .QN(n561));
   NAND2X1 U100 (.IN1(n322), .IN2(sboxw[1]), .QN(n319));
   INVX0 U101 (.INP(n1375), .ZN(n147));
   INVX0 U102 (.INP(n652), .ZN(n71));
   NAND2X1 U103 (.IN1(n211), .IN2(n228), .QN(n226));
   NAND2X1 U104 (.IN1(n563), .IN2(sboxw[25]), .QN(n560));
   INVX0 U105 (.INP(n250), .ZN(n158));
   INVX0 U106 (.INP(n563), .ZN(n74));
   NAND2X1 U107 (.IN1(n518), .IN2(n1571), .QN(n321));
   INVX0 U108 (.INP(n387), .ZN(n1545));
   NAND2X1 U109 (.IN1(n793), .IN2(n90), .QN(n562));
   NAND2X1 U110 (.IN1(n370), .IN2(n322), .QN(n352));
   NAND2X1 U111 (.IN1(n518), .IN2(n12), .QN(n476));
   NAND2X1 U112 (.IN1(n793), .IN2(n5), .QN(n717));
   INVX0 U113 (.INP(n322), .ZN(n1555));
   NAND2X1 U114 (.IN1(n611), .IN2(n563), .QN(n593));
   NOR2X0 U115 (.IN1(n79), .IN2(n87), .QN(n806));
   NAND2X1 U116 (.IN1(n387), .IN2(n12), .QN(n353));
   NAND2X1 U117 (.IN1(n206), .IN2(n28), .QN(n239));
   OA21X1 U118 (.IN1(n1552), .IN2(sboxw[1]), .IN3(n1551), .Q(n420));
   NOR2X0 U119 (.IN1(n37), .IN2(n266), .QN(n1393));
   NAND2X1 U120 (.IN1(n793), .IN2(n14), .QN(n751));
   INVX0 U121 (.INP(n628), .ZN(n64));
   INVX0 U122 (.INP(n708), .ZN(n77));
   NOR2X0 U123 (.IN1(n1560), .IN2(n1568), .QN(n531));
   NAND2X1 U124 (.IN1(n387), .IN2(n1568), .QN(n328));
   INVX0 U125 (.INP(n1048), .ZN(n120));
   NAND2X1 U126 (.IN1(n1002), .IN2(n130), .QN(n943));
   OA21X1 U127 (.IN1(n71), .IN2(sboxw[25]), .IN3(n70), .Q(n661));
   INVX0 U128 (.INP(n433), .ZN(n1558));
   INVX0 U129 (.INP(n228), .ZN(n162));
   INVX0 U130 (.INP(n568), .ZN(n59));
   INVX0 U131 (.INP(n837), .ZN(n58));
   NAND2X1 U132 (.IN1(n1164), .IN2(n13), .QN(n1091));
   NAND2X1 U133 (.IN1(n563), .IN2(n90), .QN(n752));
   NAND2X1 U134 (.IN1(n206), .IN2(n173), .QN(n1308));
   NOR2X0 U135 (.IN1(n71), .IN2(n53), .QN(n622));
   NAND2X1 U136 (.IN1(n175), .IN2(n267), .QN(n1365));
   NOR2X0 U137 (.IN1(n1568), .IN2(n1547), .QN(n365));
   INVX0 U138 (.INP(n1318), .ZN(n136));
   NAND2X1 U139 (.IN1(n628), .IN2(n14), .QN(n594));
   INVX0 U140 (.INP(n1002), .ZN(n107));
   NAND2X1 U141 (.IN1(n937), .IN2(sboxw[17]), .QN(n934));
   NOR2X0 U142 (.IN1(n1571), .IN2(n1547), .QN(n357));
   NAND2X1 U143 (.IN1(n322), .IN2(n1571), .QN(n477));
   OA21X1 U144 (.IN1(n114), .IN2(sboxw[17]), .IN3(n113), .Q(n1035));
   NOR2X0 U145 (.IN1(n87), .IN2(n66), .QN(n606));
   NAND2X1 U146 (.IN1(n1002), .IN2(n131), .QN(n1117));
   NAND2X1 U147 (.IN1(n1002), .IN2(n13), .QN(n968));
   INVX0 U148 (.INP(n599), .ZN(n50));
   NAND2X1 U149 (.IN1(n30), .IN2(n250), .QN(n224));
   NAND2X1 U150 (.IN1(n628), .IN2(n87), .QN(n569));
   NOR2X0 U151 (.IN1(n57), .IN2(n71), .QN(n817));
   NOR2X0 U152 (.IN1(n90), .IN2(n66), .QN(n598));
   NOR2X0 U153 (.IN1(n57), .IN2(n66), .QN(n896));
   NOR2X0 U154 (.IN1(n1561), .IN2(n1571), .QN(n446));
   INVX0 U155 (.INP(n582), .ZN(n82));
   INVX0 U156 (.INP(n266), .ZN(n154));
   NAND2X1 U157 (.IN1(n708), .IN2(sboxw[25]), .QN(n574));
   NOR2X0 U158 (.IN1(n100), .IN2(n109), .QN(n1267));
   NOR2X0 U159 (.IN1(n33), .IN2(n581), .QN(n716));
   INVX0 U160 (.INP(n340), .ZN(n1548));
   NAND2X1 U161 (.IN1(n1048), .IN2(sboxw[17]), .QN(n948));
   NAND2X1 U162 (.IN1(n281), .IN2(n250), .QN(n240));
   INVX0 U163 (.INP(n1166), .ZN(n104));
   INVX0 U164 (.INP(n795), .ZN(n61));
   OA21X1 U165 (.IN1(n176), .IN2(n1366), .IN3(n1329), .Q(n1471));
   NOR2X0 U166 (.IN1(n1561), .IN2(n12), .QN(n355));
   INVX0 U167 (.INP(n341), .ZN(n1563));
   NOR2X0 U168 (.IN1(n138), .IN2(n153), .QN(n290));
   NOR2X0 U169 (.IN1(n100), .IN2(n114), .QN(n1188));
   NAND2X1 U170 (.IN1(n433), .IN2(sboxw[1]), .QN(n333));
   INVX0 U171 (.INP(n520), .ZN(n1542));
   INVX0 U172 (.INP(n1208), .ZN(n101));
   INVX0 U173 (.INP(n581), .ZN(n67));
   NOR2X0 U174 (.IN1(n80), .IN2(n14), .QN(n596));
   NAND2X1 U175 (.IN1(n896), .IN2(sboxw[25]), .QN(n840));
   NOR2X0 U176 (.IN1(n80), .IN2(n90), .QN(n721));
   INVX0 U177 (.INP(n955), .ZN(n110));
   NOR2X0 U178 (.IN1(n66), .IN2(n53), .QN(n600));
   NOR2X0 U179 (.IN1(n119), .IN2(n100), .QN(n1075));
   NAND2X1 U180 (.IN1(n1267), .IN2(sboxw[17]), .QN(n1211));
   INVX0 U181 (.INP(n293), .ZN(n160));
   NOR2X0 U182 (.IN1(n143), .IN2(n159), .QN(n260));
   INVX0 U183 (.INP(n684), .ZN(n564));
   INVX0 U184 (.INP(n358), .ZN(n180));
   NAND2X1 U185 (.IN1(n1519), .IN2(sboxw[1]), .QN(n687));
   NOR2X0 U186 (.IN1(n138), .IN2(n163), .QN(n223));
   NOR2X0 U187 (.IN1(n80), .IN2(n53), .QN(n558));
   NOR2X0 U188 (.IN1(n1366), .IN2(n28), .QN(n270));
   NOR2X0 U189 (.IN1(n123), .IN2(n13), .QN(n970));
   INVX0 U190 (.INP(n1440), .ZN(n145));
   INVX0 U191 (.INP(n1316), .ZN(n168));
   INVX0 U192 (.INP(n973), .ZN(n93));
   INVX0 U193 (.INP(n956), .ZN(n125));
   INVX0 U194 (.INP(n1355), .ZN(n166));
   INVX0 U195 (.INP(n202), .ZN(n139));
   NAND2X1 U196 (.IN1(n964), .IN2(n1264), .QN(n1263));
   OR2X1 U197 (.IN1(n1571), .IN2(n39), .Q(n1));
   NOR2X0 U198 (.IN1(n35), .IN2(n179), .QN(n1139));
   NAND2X1 U199 (.IN1(n316), .IN2(n1567), .QN(n515));
   AO222X1 U200 (.IN1(n302), .IN2(n505), .IN3(n304), .IN4(n506), .IN5(n507), .IN6(n178), .
          Q(new_sboxw[3]));
   NAND2X1 U201 (.IN1(n349), .IN2(n1516), .QN(n1515));
   OA21X1 U202 (.IN1(n331), .IN2(n1546), .IN3(n393), .Q(n1537));
   INVX0 U203 (.INP(n331), .ZN(n1569));
   NAND2X1 U204 (.IN1(n590), .IN2(n893), .QN(n892));
   NOR2X0 U205 (.IN1(n931), .IN2(n1048), .QN(n1046));
   INVX0 U206 (.INP(n1047), .ZN(n124));
   OA21X1 U207 (.IN1(n316), .IN2(n322), .IN3(n1567), .Q(n532));
   NOR2X0 U208 (.IN1(n316), .IN2(n433), .QN(n431));
   INVX0 U209 (.INP(n432), .ZN(n1562));
   OA222X1 U210 (.IN1(n129), .IN2(n123), .IN3(n131), .IN4(n108), .IN5(n107), .IN6(n32), .Q(
          n1236));
   NAND2X1 U211 (.IN1(n128), .IN2(n115), .QN(n1237));
   OA21X1 U212 (.IN1(n131), .IN2(n111), .IN3(n1038), .Q(n1272));
   AO22X1 U213 (.IN1(n922), .IN2(n1195), .IN3(n988), .IN4(n1196), .Q(n1194));
   OAI222X1 U214 (.IN1(n108), .IN2(n31), .IN3(n1090), .IN4(n946), .IN5(n118), .IN6(n13), .
          QN(n1089));
   NOR2X0 U215 (.IN1(n557), .IN2(n708), .QN(n706));
   INVX0 U216 (.INP(n707), .ZN(n81));
   NOR2X0 U217 (.IN1(n1166), .IN2(n1006), .QN(n1221));
   INVX0 U218 (.INP(n572), .ZN(n88));
   NAND2X1 U219 (.IN1(n1186), .IN2(n938), .QN(n1106));
   NOR2X0 U220 (.IN1(n520), .IN2(n391), .QN(n697));
   NAND2X1 U221 (.IN1(n557), .IN2(n86), .QN(n790));
   NOR2X0 U222 (.IN1(n33), .IN2(n49), .QN(n871));
   NOR2X0 U223 (.IN1(n938), .IN2(n92), .QN(n1242));
   OA21X1 U224 (.IN1(n1011), .IN2(n111), .IN3(n121), .Q(n1205));
   NAND2X1 U225 (.IN1(n1566), .IN2(n1553), .QN(n1134));
   NAND2X1 U226 (.IN1(n938), .IN2(n937), .QN(n1099));
   NAND3X0 U227 (.IN1(n957), .IN2(n128), .IN3(n955), .QN(n1101));
   OA21X1 U228 (.IN1(n396), .IN2(n1549), .IN3(n1559), .Q(n681));
   OA21X1 U229 (.IN1(n1569), .IN2(n1549), .IN3(n423), .Q(n1524));
   NAND2X1 U230 (.IN1(n938), .IN2(n115), .QN(n1115));
   OA21X1 U231 (.IN1(n572), .IN2(n65), .IN3(n634), .Q(n914));
   NOR2X0 U232 (.IN1(n370), .IN2(n339), .QN(n537));
   NAND2X1 U233 (.IN1(n817), .IN2(n86), .QN(n898));
   INVX0 U234 (.INP(n1011), .ZN(n130));
   NAND2X1 U235 (.IN1(n130), .IN2(n128), .QN(n1016));
   AO222X1 U236 (.IN1(n543), .IN2(n544), .IN3(n545), .IN4(n546), .IN5(n547), .IN6(n48), .Q(
          new_sboxw[31]));
   NAND2X1 U237 (.IN1(n601), .IN2(n602), .QN(n544));
   NOR2X0 U238 (.IN1(n1566), .IN2(n1552), .QN(n518));
   NOR2X0 U239 (.IN1(n1553), .IN2(n1564), .QN(n411));
   NAND2X1 U240 (.IN1(n1), .IN2(n349), .QN(n348));
   NAND2X1 U241 (.IN1(n35), .IN2(n1553), .QN(n500));
   INVX0 U242 (.INP(n1300), .ZN(n146));
   NOR2X0 U243 (.IN1(n155), .IN2(n167), .QN(n244));
   NAND2X1 U244 (.IN1(n158), .IN2(n146), .QN(n1469));
   NAND2X1 U245 (.IN1(n540), .IN2(n35), .QN(n491));
   OA21X1 U246 (.IN1(n557), .IN2(n563), .IN3(n86), .Q(n807));
   OR2X1 U247 (.IN1(n90), .IN2(n46), .Q(n2));
   NAND2X1 U248 (.IN1(n391), .IN2(n39), .QN(n389));
   NOR2X0 U249 (.IN1(n153), .IN2(n172), .QN(n206));
   INVX0 U250 (.INP(n241), .ZN(n153));
   INVX0 U251 (.INP(n262), .ZN(n151));
   NAND2X0 U252 (.IN1(n35), .IN2(n322), .QN(n484));
   OA21X1 U253 (.IN1(n88), .IN2(n68), .IN3(n664), .Q(n901));
   NOR2X0 U254 (.IN1(n1186), .IN2(n937), .QN(n1253));
   NOR2X0 U255 (.IN1(n795), .IN2(n632), .QN(n850));
   NOR2X0 U256 (.IN1(n115), .IN2(n126), .QN(n1026));
   OA21X1 U257 (.IN1(n637), .IN2(n68), .IN3(n78), .Q(n834));
   AO222X1 U258 (.IN1(n1288), .IN2(n1289), .IN3(n1290), .IN4(n1291), .IN5(n1292), .IN6(
          n134), .Q(new_sboxw[15]));
   NAND2X1 U259 (.IN1(n1326), .IN2(n1327), .QN(n1289));
   AO22X1 U260 (.IN1(n990), .IN2(n1157), .IN3(n988), .IN4(n1158), .Q(n1156));
   NAND2X1 U261 (.IN1(n331), .IN2(n391), .QN(n346));
   NOR2X0 U262 (.IN1(n148), .IN2(n172), .QN(n1375));
   INVX0 U263 (.INP(n557), .ZN(n68));
   NOR2X0 U264 (.IN1(n72), .IN2(n83), .QN(n652));
   NAND2X1 U265 (.IN1(n85), .IN2(n72), .QN(n866));
   NAND2X1 U266 (.IN1(n975), .IN2(n976), .QN(n918));
   NOR2X0 U267 (.IN1(n37), .IN2(n135), .QN(n222));
   NOR2X0 U268 (.IN1(n85), .IN2(n71), .QN(n793));
   NOR2X0 U269 (.IN1(n172), .IN2(n159), .QN(n250));
   INVX0 U270 (.INP(n245), .ZN(n159));
   INVX0 U271 (.INP(n931), .ZN(n111));
   NOR2X0 U272 (.IN1(n76), .IN2(n85), .QN(n563));
   NAND2X0 U273 (.IN1(n33), .IN2(n563), .QN(n759));
   NAND2X1 U274 (.IN1(n391), .IN2(n6), .QN(n434));
   OA21X1 U275 (.IN1(n1555), .IN2(n331), .IN3(n321), .Q(n368));
   INVX0 U276 (.INP(n316), .ZN(n1549));
   NAND2X1 U277 (.IN1(n1375), .IN2(n177), .QN(n1305));
   OA21X1 U278 (.IN1(n158), .IN2(n204), .IN3(n1305), .Q(n1333));
   INVX0 U279 (.INP(n1372), .ZN(n170));
   NOR2X0 U280 (.IN1(n1566), .IN2(n1547), .QN(n387));
   INVX0 U281 (.INP(n447), .ZN(n1547));
   NAND2X1 U282 (.IN1(n396), .IN2(n387), .QN(n478));
   NOR2X0 U283 (.IN1(n228), .IN2(n249), .QN(n1315));
   OA21X1 U284 (.IN1(n74), .IN2(n572), .IN3(n562), .Q(n609));
   OA21X1 U285 (.IN1(n1571), .IN2(n480), .IN3(n1551), .Q(n479));
   NOR2X0 U286 (.IN1(n386), .IN2(n387), .QN(n384));
   INVX0 U287 (.INP(n540), .ZN(n1546));
   NOR2X0 U288 (.IN1(n985), .IN2(n954), .QN(n1183));
   NOR2X0 U289 (.IN1(n433), .IN2(n540), .QN(n339));
   INVX0 U290 (.INP(n249), .ZN(n150));
   OA21X1 U291 (.IN1(n177), .IN2(n265), .IN3(n147), .Q(n1421));
   NOR2X0 U292 (.IN1(n1557), .IN2(n1566), .QN(n322));
   NAND2X1 U293 (.IN1(n37), .IN2(n250), .QN(n1425));
   INVX0 U294 (.INP(n590), .ZN(n80));
   INVX0 U295 (.INP(n627), .ZN(n79));
   NAND2X1 U296 (.IN1(n563), .IN2(n4), .QN(n664));
   INVX0 U297 (.INP(n334), .ZN(n1565));
   NAND2X1 U298 (.IN1(n331), .IN2(n1566), .QN(n392));
   INVX0 U299 (.INP(n1470), .ZN(n157));
   NAND2X1 U300 (.IN1(n245), .IN2(n174), .QN(n1387));
   NAND2X1 U301 (.IN1(n37), .IN2(n155), .QN(n1441));
   INVX0 U302 (.INP(n964), .ZN(n123));
   INVX0 U303 (.INP(n1001), .ZN(n122));
   INVX0 U304 (.INP(n722), .ZN(n66));
   NOR2X0 U305 (.IN1(n708), .IN2(n815), .QN(n580));
   INVX0 U306 (.INP(n359), .ZN(n182));
   NAND2X1 U307 (.IN1(n37), .IN2(n249), .QN(n1432));
   NAND2X1 U308 (.IN1(n1489), .IN2(n1490), .QN(n1480));
   NOR2X0 U309 (.IN1(n85), .IN2(n66), .QN(n628));
   OA21X1 U310 (.IN1(n90), .IN2(n755), .IN3(n70), .Q(n754));
   NOR2X0 U311 (.IN1(n85), .IN2(n80), .QN(n708));
   INVX0 U312 (.INP(n632), .ZN(n76));
   NAND2X1 U313 (.IN1(n572), .IN2(n632), .QN(n587));
   INVX0 U314 (.INP(n815), .ZN(n65));
   NAND2X1 U315 (.IN1(n300), .IN2(n37), .QN(n1422));
   INVX0 U316 (.INP(n349), .ZN(n1561));
   INVX0 U317 (.INP(n386), .ZN(n1560));
   NOR2X0 U318 (.IN1(n518), .IN2(n541), .QN(n679));
   NOR2X0 U319 (.IN1(n119), .IN2(n128), .QN(n937));
   NOR2X0 U320 (.IN1(n1375), .IN2(n1470), .QN(n212));
   NAND2X1 U321 (.IN1(n637), .IN2(n628), .QN(n753));
   NOR2X0 U322 (.IN1(n639), .IN2(n11), .QN(n715));
   NAND2X1 U323 (.IN1(n582), .IN2(n72), .QN(n639));
   NAND2X1 U324 (.IN1(n774), .IN2(n750), .QN(n582));
   NOR2X0 U325 (.IN1(n128), .IN2(n123), .QN(n1048));
   INVX0 U326 (.INP(n1062), .ZN(n109));
   INVX0 U327 (.INP(n1186), .ZN(n108));
   NOR2X0 U328 (.IN1(n793), .IN2(n816), .QN(n832));
   INVX0 U329 (.INP(n575), .ZN(n84));
   NOR2X0 U330 (.IN1(n1566), .IN2(n1561), .QN(n433));
   NAND2X1 U331 (.IN1(n632), .IN2(n5), .QN(n709));
   INVX0 U332 (.INP(n197), .ZN(n171));
   NOR2X0 U333 (.IN1(n163), .IN2(n172), .QN(n228));
   INVX0 U334 (.INP(n242), .ZN(n163));
   INVX0 U335 (.INP(n391), .ZN(n1557));
   INVX0 U336 (.INP(n715), .ZN(n60));
   NAND2X1 U337 (.IN1(n32), .IN2(n964), .QN(n963));
   NAND2X1 U338 (.IN1(n1011), .IN2(n1002), .QN(n1093));
   OA21X1 U339 (.IN1(n133), .IN2(n1095), .IN3(n113), .Q(n1094));
   NAND2X1 U340 (.IN1(n637), .IN2(n563), .QN(n720));
   NOR2X0 U341 (.IN1(n85), .IN2(n11), .QN(n568));
   NOR2X0 U342 (.IN1(n59), .IN2(n83), .QN(n837));
   OA21X1 U343 (.IN1(n211), .IN2(n157), .IN3(n1371), .Q(n1491));
   NAND2X1 U344 (.IN1(n250), .IN2(n3), .QN(n214));
   NOR2X0 U345 (.IN1(n46), .IN2(n51), .QN(n599));
   INVX0 U346 (.INP(n204), .ZN(n175));
   INVX0 U347 (.INP(n816), .ZN(n75));
   NOR2X0 U348 (.IN1(n92), .IN2(n45), .QN(n924));
   NAND2X1 U349 (.IN1(n572), .IN2(n85), .QN(n633));
   NAND2X1 U350 (.IN1(n387), .IN2(n39), .QN(n698));
   NAND2X1 U351 (.IN1(n1011), .IN2(n937), .QN(n1060));
   NAND2X1 U352 (.IN1(n628), .IN2(n46), .QN(n851));
   NAND2X1 U353 (.IN1(n250), .IN2(n177), .QN(n208));
   NAND2X1 U354 (.IN1(n341), .IN2(n1553), .QN(n398));
   NAND2X1 U355 (.IN1(n499), .IN2(n475), .QN(n341));
   NAND2X1 U356 (.IN1(n396), .IN2(n322), .QN(n445));
   OAI221X1 U357 (.IN1(n120), .IN2(n946), .IN3(n117), .IN4(n1011), .IN5(n1091), .QN(n1277)
          );
   NOR2X0 U358 (.IN1(n1164), .IN2(n1187), .QN(n1203));
   INVX0 U359 (.INP(n201), .ZN(n173));
   NAND2X1 U360 (.IN1(n173), .IN2(n172), .QN(n267));
   INVX0 U361 (.INP(n1349), .ZN(n161));
   INVX0 U362 (.INP(n541), .ZN(n1556));
   OA222X1 U363 (.IN1(n946), .IN2(n113), .IN3(n133), .IN4(n947), .IN5(n938), .IN6(n111), .
          Q(n945));
   INVX0 U364 (.INP(n949), .ZN(n127));
   NOR2X0 U365 (.IN1(n1300), .IN2(n228), .QN(n1386));
   NAND2X1 U366 (.IN1(n1002), .IN2(n44), .QN(n1222));
   NAND3X0 U367 (.IN1(n1568), .IN2(n1547), .IN3(n366), .QN(n688));
   INVX0 U368 (.INP(n440), .ZN(n1541));
   INVX0 U369 (.INP(n1006), .ZN(n119));
   NOR2X0 U370 (.IN1(n56), .IN2(n637), .QN(n646));
   NAND2X1 U371 (.IN1(n433), .IN2(n40), .QN(n326));
   OA21X1 U372 (.IN1(n1553), .IN2(n323), .IN3(n326), .Q(n324));
   NAND2X1 U373 (.IN1(n815), .IN2(n33), .QN(n766));
   NAND2X1 U374 (.IN1(n85), .IN2(n83), .QN(n573));
   NOR2X0 U375 (.IN1(n44), .IN2(n94), .QN(n973));
   NOR2X0 U376 (.IN1(n242), .IN2(n241), .QN(n266));
   NOR2X0 U377 (.IN1(n99), .IN2(n1011), .QN(n1020));
   NAND2X1 U378 (.IN1(n228), .IN2(n43), .QN(n194));
   OA21X1 U379 (.IN1(n155), .IN2(n143), .IN3(n194), .Q(n1306));
   NOR2X0 U380 (.IN1(n349), .IN2(n447), .QN(n340));
   NAND2X1 U381 (.IN1(n87), .IN2(n85), .QN(n642));
   NOR2X0 U382 (.IN1(n128), .IN2(n115), .QN(n1166));
   NOR2X0 U383 (.IN1(n85), .IN2(n72), .QN(n795));
   OA21X1 U384 (.IN1(n72), .IN2(n57), .IN3(n567), .Q(n565));
   NAND2X1 U385 (.IN1(n128), .IN2(n126), .QN(n947));
   INVX0 U386 (.INP(n1187), .ZN(n118));
   NAND2X1 U387 (.IN1(n1566), .IN2(n1564), .QN(n332));
   INVX0 U388 (.INP(n1055), .ZN(n103));
   NAND2X1 U389 (.IN1(n33), .IN2(n72), .QN(n775));
   INVX0 U390 (.INP(n607), .ZN(n57));
   NAND2X1 U391 (.IN1(n1568), .IN2(n1566), .QN(n401));
   NOR2X0 U392 (.IN1(n1566), .IN2(n1553), .QN(n520));
   NAND2X1 U393 (.IN1(n1547), .IN2(n1566), .QN(n676));
   NAND2X1 U394 (.IN1(n29), .IN2(n1349), .QN(n1371));
   NOR2X0 U395 (.IN1(n590), .IN2(n722), .QN(n581));
   NAND2X1 U396 (.IN1(n153), .IN2(n172), .QN(n1488));
   NOR2X0 U397 (.IN1(n102), .IN2(n126), .QN(n1208));
   INVX0 U398 (.INP(n942), .ZN(n102));
   NAND2X1 U399 (.IN1(n1114), .IN2(n1090), .QN(n956));
   NAND2X1 U400 (.IN1(n956), .IN2(n115), .QN(n1013));
   NOR2X0 U401 (.IN1(n964), .IN2(n1062), .QN(n955));
   NAND2X1 U402 (.IN1(n66), .IN2(n85), .QN(n829));
   NOR2X0 U403 (.IN1(n92), .IN2(n91), .QN(n917));
   NAND2X1 U404 (.IN1(n109), .IN2(n128), .QN(n1200));
   NAND2X1 U405 (.IN1(n1048), .IN2(n45), .QN(n941));
   NOR2X0 U406 (.IN1(n177), .IN2(n163), .QN(n293));
   NAND2X1 U407 (.IN1(n627), .IN2(n14), .QN(n577));
   NAND2X1 U408 (.IN1(n29), .IN2(n241), .QN(n1331));
   NAND2X1 U409 (.IN1(n600), .IN2(n46), .QN(n584));
   NAND2X1 U410 (.IN1(n386), .IN2(n12), .QN(n336));
   NAND2X1 U411 (.IN1(n173), .IN2(n43), .QN(n1307));
   NAND2X1 U412 (.IN1(n130), .IN2(n45), .QN(n940));
   NAND2X1 U413 (.IN1(n1001), .IN2(n13), .QN(n951));
   NAND2X1 U414 (.IN1(n286), .IN2(n241), .QN(n1366));
   NAND2X1 U415 (.IN1(n359), .IN2(n39), .QN(n343));
   NAND3X0 U416 (.IN1(n41), .IN2(n154), .IN3(n286), .QN(n1463));
   INVX0 U417 (.INP(n739), .ZN(n53));
   NOR2X0 U418 (.IN1(n1048), .IN2(n1186), .QN(n954));
   NOR2X0 U419 (.IN1(n155), .IN2(n172), .QN(n1440));
   OA21X1 U420 (.IN1(n115), .IN2(n100), .IN3(n941), .Q(n939));
   NAND2X1 U421 (.IN1(n300), .IN2(n204), .QN(n1484));
   NAND2X1 U422 (.IN1(n217), .IN2(n169), .QN(n1316));
   INVX0 U423 (.INP(n1354), .ZN(n164));
   NAND2X1 U424 (.IN1(n632), .IN2(n46), .QN(n630));
   INVX0 U425 (.INP(n1348), .ZN(n165));
   NAND2X1 U426 (.IN1(n1006), .IN2(n44), .QN(n1004));
   NAND2X1 U427 (.IN1(n974), .IN2(n44), .QN(n958));
   INVX0 U428 (.INP(n637), .ZN(n87));
   NOR2X0 U429 (.IN1(n49), .IN2(n11), .QN(n548));
   INVX0 U430 (.INP(n396), .ZN(n1568));
   NOR2X0 U431 (.IN1(n179), .IN2(n40), .QN(n309));
   NOR2X0 U432 (.IN1(n167), .IN2(n172), .QN(n1355));
   NAND2X1 U433 (.IN1(n172), .IN2(n167), .QN(n237));
   NOR2X0 U434 (.IN1(n140), .IN2(n167), .QN(n202));
   NOR2X0 U435 (.IN1(n49), .IN2(n48), .QN(n543));
   NOR2X0 U436 (.IN1(n179), .IN2(n178), .QN(n302));
   NAND2X1 U437 (.IN1(n1568), .IN2(n40), .QN(n325));
   INVX0 U438 (.INP(n299), .ZN(n169));
   NOR2X0 U439 (.IN1(n135), .IN2(n43), .QN(n190));
   NOR2X0 U440 (.IN1(n134), .IN2(n135), .QN(n1288));
   INVX0 U441 (.INP(n271), .ZN(n140));
   INVX0 U442 (.INP(n229), .ZN(n138));
   AO22X1 U443 (.IN1(n1256), .IN2(n92), .IN3(sboxw[22]), .IN4(n1257), .Q(n1255));
   INVX0 U444 (.INP(n21), .ZN(n133));
   NAND2X1 U445 (.IN1(n1282), .IN2(n132), .QN(n1264));
   NAND2X1 U446 (.IN1(n1188), .IN2(n21), .QN(n1259));
   INVX0 U447 (.INP(n1020), .ZN(n98));
   OA21X1 U448 (.IN1(n955), .IN2(n1016), .IN3(n1204), .Q(n1265));
   AO222X1 U449 (.IN1(n919), .IN2(n1039), .IN3(n1040), .IN4(n91), .IN5(n917), .IN6(n1041)
          , .Q(new_sboxw[21]));
   AO22X1 U450 (.IN1(n1050), .IN2(n92), .IN3(sboxw[22]), .IN4(n1051), .Q(n1040));
   AO221X1 U451 (.IN1(n981), .IN2(n1052), .IN3(n10), .IN4(n1053), .IN5(n1054), .Q(n1051)
          );
   NAND2X1 U452 (.IN1(n997), .IN2(n998), .QN(n994));
   NAND2X1 U453 (.IN1(n1027), .IN2(n1028), .QN(n1018));
   AO22X1 U454 (.IN1(sboxw[7]), .IN2(n1120), .IN3(n1121), .IN4(n178), .Q(new_sboxw[1]));
   NAND2X1 U455 (.IN1(n1534), .IN2(n1570), .QN(n1516));
   NAND2X1 U456 (.IN1(n542), .IN2(n15), .QN(n1511));
   AO22X1 U457 (.IN1(sboxw[7]), .IN2(n1506), .IN3(n1507), .IN4(n178), .Q(new_sboxw[0]));
   AOI222X1 U458 (.IN1(n8), .IN2(n1513), .IN3(n1514), .IN4(n40), .IN5(n460), .IN6(n39), .
          QN(n1512));
   OA21X1 U459 (.IN1(n340), .IN2(n401), .IN3(n680), .Q(n1517));
   AO222X1 U460 (.IN1(n304), .IN2(n424), .IN3(n425), .IN4(n178), .IN5(n302), .IN6(n426), .
          Q(new_sboxw[5]));
   NAND2X1 U461 (.IN1(n1186), .IN2(n132), .QN(n1214));
   AO22X1 U462 (.IN1(n371), .IN2(n178), .IN3(sboxw[7]), .IN4(n372), .Q(new_sboxw[6]));
   NAND2X1 U463 (.IN1(n412), .IN2(n413), .QN(n403));
   OA21X1 U464 (.IN1(n17), .IN2(n396), .IN3(sboxw[3]), .Q(n415));
   NAND2X1 U465 (.IN1(n23), .IN2(n132), .QN(n1077));
   NOR2X0 U466 (.IN1(sboxw[3]), .IN2(n323), .QN(n1535));
   NOR2X0 U467 (.IN1(n12), .IN2(n15), .QN(n331));
   NAND2X1 U468 (.IN1(n407), .IN2(n408), .QN(n406));
   NAND2X1 U469 (.IN1(n911), .IN2(n89), .QN(n893));
   NAND2X1 U470 (.IN1(n817), .IN2(n24), .QN(n888));
   INVX0 U471 (.INP(n646), .ZN(n55));
   OA21X1 U472 (.IN1(n581), .IN2(n642), .IN3(n833), .Q(n894));
   OA21X1 U473 (.IN1(n1070), .IN2(n100), .IN3(n97), .Q(n1063));
   OA21X1 U474 (.IN1(n985), .IN2(n126), .IN3(n32), .Q(n1070));
   NOR2X0 U475 (.IN1(sboxw[19]), .IN2(n100), .QN(n1283));
   AOI222X1 U476 (.IN1(n8), .IN2(n1523), .IN3(n440), .IN4(n1569), .IN5(n460), .IN6(n1570)
          , .QN(n1522));
   NAND2X1 U477 (.IN1(n542), .IN2(n1567), .QN(n1521));
   OA21X1 U478 (.IN1(n455), .IN2(n323), .IN3(n184), .Q(n448));
   OA21X1 U479 (.IN1(n370), .IN2(n1564), .IN3(n1), .Q(n455));
   NOR2X0 U480 (.IN1(n39), .IN2(n1556), .QN(n530));
   NAND2X1 U481 (.IN1(n17), .IN2(n1570), .QN(n462));
   NAND2X1 U482 (.IN1(n1251), .IN2(n1252), .QN(n1238));
   AO22X1 U483 (.IN1(n990), .IN2(n1105), .IN3(n985), .IN4(n996), .Q(n1104));
   AO221X1 U484 (.IN1(n988), .IN2(n1102), .IN3(sboxw[22]), .IN4(n1103), .IN5(n1104), .Q(
          n1080));
   NAND3X0 U485 (.IN1(n957), .IN2(n110), .IN3(n942), .QN(n1268));
   NOR2X0 U486 (.IN1(n1088), .IN2(n1089), .QN(n1087));
   AO222X1 U487 (.IN1(n302), .IN2(n665), .IN3(n304), .IN4(n666), .IN5(n667), .IN6(n178), .
          Q(new_sboxw[2]));
   NOR2X0 U488 (.IN1(n1011), .IN2(n955), .QN(n1281));
   NOR2X0 U489 (.IN1(n14), .IN2(n24), .QN(n572));
   AO22X1 U490 (.IN1(n612), .IN2(n48), .IN3(sboxw[31]), .IN4(n613), .Q(new_sboxw[30]));
   NAND2X1 U491 (.IN1(n648), .IN2(n649), .QN(n647));
   NAND2X1 U492 (.IN1(n540), .IN2(n1570), .QN(n690));
   OA21X1 U493 (.IN1(n1567), .IN2(n1558), .IN3(n368), .Q(n691));
   AO22X1 U494 (.IN1(sboxw[31]), .IN2(n852), .IN3(n853), .IN4(n48), .Q(new_sboxw[25]));
   NAND2X1 U495 (.IN1(n35), .IN2(sboxw[3]), .QN(n416));
   NAND2X1 U496 (.IN1(n26), .IN2(n89), .QN(n737));
   NOR2X0 U497 (.IN1(n721), .IN2(n597), .QN(n738));
   NAND2X1 U498 (.IN1(n382), .IN2(n383), .QN(n379));
   NOR2X0 U499 (.IN1(n597), .IN2(n793), .QN(n803));
   NOR2X0 U500 (.IN1(n46), .IN2(n75), .QN(n805));
   NAND2X1 U501 (.IN1(n653), .IN2(n654), .QN(n644));
   OA21X1 U502 (.IN1(n26), .IN2(n637), .IN3(sboxw[27]), .Q(n656));
   NOR2X0 U503 (.IN1(sboxw[27]), .IN2(n57), .QN(n912));
   OA221X1 U504 (.IN1(n957), .IN2(n108), .IN3(n21), .IN4(n999), .IN5(n1000), .Q(n998));
   OA21X1 U505 (.IN1(n109), .IN2(n131), .IN3(n982), .Q(n1074));
   OA21X1 U506 (.IN1(n107), .IN2(n32), .IN3(n1060), .Q(n1076));
   OA21X1 U507 (.IN1(n730), .IN2(n57), .IN3(n54), .Q(n723));
   OA21X1 U508 (.IN1(n611), .IN2(n83), .IN3(n2), .Q(n730));
   NAND2X1 U509 (.IN1(n22), .IN2(sboxw[19]), .QN(n1012));
   OA21X1 U510 (.IN1(n21), .IN2(n1012), .IN3(n113), .Q(n1065));
   NOR2X0 U511 (.IN1(n44), .IN2(n21), .QN(n1011));
   NAND2X1 U512 (.IN1(n1022), .IN2(n1023), .QN(n1021));
   NAND2X1 U513 (.IN1(n623), .IN2(n624), .QN(n620));
   INVX0 U514 (.INP(n17), .ZN(n1553));
   AO22X1 U515 (.IN1(n740), .IN2(n48), .IN3(sboxw[31]), .IN4(n741), .Q(new_sboxw[28]));
   OA21X1 U516 (.IN1(n86), .IN2(n77), .IN3(n609), .Q(n844));
   NAND2X1 U517 (.IN1(n815), .IN2(n89), .QN(n843));
   INVX0 U518 (.INP(n18), .ZN(n177));
   NOR2X0 U519 (.IN1(sboxw[11]), .IN2(n173), .QN(n294));
   NAND2X1 U520 (.IN1(n1367), .IN2(n1368), .QN(n1359));
   OA21X1 U521 (.IN1(n20), .IN2(n27), .IN3(sboxw[11]), .Q(n1370));
   NOR2X0 U522 (.IN1(n396), .IN2(n340), .QN(n1533));
   INVX0 U523 (.INP(n20), .ZN(n155));
   NOR2X0 U524 (.IN1(n148), .IN2(n19), .QN(n1300));
   NOR2X0 U525 (.IN1(n149), .IN2(n1375), .QN(n1466));
   NOR2X0 U526 (.IN1(n1467), .IN2(n1468), .QN(n1465));
   AO22X1 U527 (.IN1(n375), .IN2(n490), .IN3(n370), .IN4(n381), .Q(n489));
   AOI222X1 U528 (.IN1(n8), .IN2(n364), .IN3(n365), .IN4(n40), .IN5(n355), .IN6(n366), .QN(
          n360));
   OA21X1 U529 (.IN1(n1403), .IN2(n143), .IN3(n142), .Q(n1396));
   OA21X1 U530 (.IN1(n281), .IN2(n167), .IN3(n3), .Q(n1403));
   NOR2X0 U531 (.IN1(n473), .IN2(n474), .QN(n472));
   AO221X1 U532 (.IN1(n249), .IN2(n176), .IN3(n1300), .IN4(n42), .IN5(n1353), .Q(n1340));
   OA21X1 U533 (.IN1(n1547), .IN2(n1569), .IN3(n367), .Q(n459));
   OA21X1 U534 (.IN1(n1545), .IN2(n1), .IN3(n445), .Q(n461));
   OA21X1 U535 (.IN1(n266), .IN2(n267), .IN3(n268), .Q(n263));
   NOR2X0 U536 (.IN1(n155), .IN2(sboxw[11]), .QN(n241));
   OR2X1 U537 (.IN1(n177), .IN2(n42), .Q(n3));
   NAND2X1 U538 (.IN1(n37), .IN2(sboxw[11]), .QN(n236));
   NAND2X1 U539 (.IN1(n20), .IN2(n176), .QN(n1409));
   NOR2X0 U540 (.IN1(n293), .IN2(n149), .QN(n1410));
   INVX0 U541 (.INP(n23), .ZN(n115));
   NOR2X0 U542 (.IN1(n748), .IN2(n749), .QN(n747));
   NOR2X0 U543 (.IN1(n1474), .IN2(n1475), .QN(n1473));
   OAI221X1 U544 (.IN1(n1315), .IN2(n281), .IN3(n161), .IN4(n30), .IN5(n214), .QN(n1474)
          );
   NAND2X1 U545 (.IN1(n1148), .IN2(n1149), .QN(n1135));
   NOR2X0 U546 (.IN1(n540), .IN2(n322), .QN(n1150));
   NOR2X0 U547 (.IN1(n611), .IN2(n580), .QN(n812));
   NOR2X0 U548 (.IN1(n44), .IN2(n118), .QN(n1176));
   INVX0 U549 (.INP(n26), .ZN(n72));
   NOR2X0 U550 (.IN1(n71), .IN2(n25), .QN(n557));
   NOR2X0 U551 (.IN1(n1349), .IN2(n206), .QN(n1347));
   NAND2X1 U552 (.IN1(n1345), .IN2(n1346), .QN(n1343));
   NOR2X0 U553 (.IN1(sboxw[11]), .IN2(n20), .QN(n245));
   NOR2X0 U554 (.IN1(n114), .IN2(n22), .QN(n931));
   INVX0 U555 (.INP(n16), .ZN(n1566));
   OA21X1 U556 (.IN1(n572), .IN2(n910), .IN3(n11), .Q(n908));
   NOR2X0 U557 (.IN1(n637), .IN2(n581), .QN(n910));
   NAND2X1 U558 (.IN1(n2), .IN2(n590), .QN(n589));
   INVX0 U559 (.INP(n25), .ZN(n85));
   NOR2X0 U560 (.IN1(n1552), .IN2(n16), .QN(n316));
   NOR2X0 U561 (.IN1(n1553), .IN2(sboxw[3]), .QN(n447));
   NOR2X0 U562 (.IN1(n153), .IN2(n19), .QN(n249));
   OA21X1 U563 (.IN1(n153), .IN2(n175), .IN3(n1334), .Q(n1407));
   OA21X1 U564 (.IN1(n152), .IN2(n3), .IN3(n224), .Q(n1408));
   AO222X1 U565 (.IN1(n1288), .IN2(n1476), .IN3(n1290), .IN4(n1477), .IN5(n1478), .IN6(
          n134), .Q(new_sboxw[10]));
   NOR2X0 U566 (.IN1(n1547), .IN2(n16), .QN(n540));
   NAND2X1 U567 (.IN1(n518), .IN2(n15), .QN(n409));
   OA21X1 U568 (.IN1(n204), .IN2(n159), .IN3(n1325), .Q(n1417));
   NOR2X0 U569 (.IN1(n1419), .IN2(n1420), .QN(n1418));
   OA21X1 U570 (.IN1(n15), .IN2(n397), .IN3(n1551), .Q(n450));
   NOR2X0 U571 (.IN1(n83), .IN2(n26), .QN(n590));
   NOR2X0 U572 (.IN1(n80), .IN2(n25), .QN(n627));
   OA21X1 U573 (.IN1(n18), .IN2(n166), .IN3(n147), .Q(n1398));
   OA21X1 U574 (.IN1(n66), .IN2(n88), .IN3(n608), .Q(n734));
   OA21X1 U575 (.IN1(n64), .IN2(n2), .IN3(n720), .Q(n736));
   NOR2X0 U576 (.IN1(n159), .IN2(n19), .QN(n1470));
   NAND2X1 U577 (.IN1(n249), .IN2(n176), .QN(n1498));
   OA21X1 U578 (.IN1(n211), .IN2(n162), .IN3(n1333), .Q(n1499));
   NAND2X1 U579 (.IN1(n246), .IN2(n247), .QN(n218));
   NOR2X0 U580 (.IN1(n249), .IN2(n250), .QN(n248));
   NAND2X1 U581 (.IN1(n37), .IN2(n1349), .QN(n1456));
   NOR2X0 U582 (.IN1(n126), .IN2(n23), .QN(n964));
   NOR2X0 U583 (.IN1(n123), .IN2(n22), .QN(n1001));
   AOI222X1 U584 (.IN1(n1300), .IN2(n41), .IN3(n223), .IN4(n175), .IN5(n9), .IN6(n1301), .
          QN(n1299));
   NOR2X0 U585 (.IN1(n66), .IN2(n25), .QN(n815));
   NAND2X1 U586 (.IN1(n880), .IN2(n881), .QN(n867));
   NOR2X0 U587 (.IN1(n815), .IN2(n563), .QN(n882));
   NAND2X1 U588 (.IN1(n793), .IN2(n24), .QN(n650));
   OA21X1 U589 (.IN1(n24), .IN2(n638), .IN3(n70), .Q(n725));
   NAND2X1 U590 (.IN1(n1375), .IN2(n18), .QN(n1364));
   NAND2X1 U591 (.IN1(n1365), .IN2(n155), .QN(n1362));
   NOR2X0 U592 (.IN1(sboxw[27]), .IN2(n26), .QN(n632));
   NOR2X0 U593 (.IN1(n1564), .IN2(n17), .QN(n349));
   NOR2X0 U594 (.IN1(n1561), .IN2(n16), .QN(n386));
   INVX0 U595 (.INP(n22), .ZN(n128));
   NAND2X1 U596 (.IN1(sboxw[27]), .IN2(n85), .QN(n750));
   NOR2X0 U597 (.IN1(n109), .IN2(n22), .QN(n1186));
   NOR2X0 U598 (.IN1(n627), .IN2(n628), .QN(n625));
   INVX0 U599 (.INP(n600), .ZN(n52));
   NOR2X0 U600 (.IN1(n167), .IN2(n20), .QN(n242));
   NOR2X0 U601 (.IN1(sboxw[3]), .IN2(n17), .QN(n391));
   NAND2X1 U602 (.IN1(n33), .IN2(sboxw[27]), .QN(n657));
   OA222X1 U603 (.IN1(n211), .IN2(n146), .IN3(n1504), .IN4(n42), .IN5(n176), .IN6(n265), .
          Q(n1503));
   NOR2X0 U604 (.IN1(n1440), .IN2(n245), .QN(n1504));
   NAND3X0 U605 (.IN1(n23), .IN2(n956), .IN3(n957), .QN(n950));
   NOR2X0 U606 (.IN1(n76), .IN2(n25), .QN(n816));
   NAND3X0 U607 (.IN1(n129), .IN2(n126), .IN3(n942), .QN(n927));
   INVX0 U608 (.INP(sboxw[22]), .ZN(n92));
   INVX0 U609 (.INP(n42), .ZN(n41));
   NAND2X1 U610 (.IN1(sboxw[3]), .IN2(n1566), .QN(n475));
   NOR2X0 U611 (.IN1(n163), .IN2(n19), .QN(n1349));
   NOR2X0 U612 (.IN1(n1557), .IN2(n16), .QN(n541));
   NOR2X0 U613 (.IN1(n92), .IN2(n10), .QN(n922));
   NOR2X0 U614 (.IN1(n27), .IN2(n266), .QN(n292));
   NOR2X0 U615 (.IN1(n119), .IN2(n22), .QN(n1187));
   NOR2X0 U616 (.IN1(n25), .IN2(n11), .QN(n607));
   NAND2X1 U617 (.IN1(n281), .IN2(n19), .QN(n1453));
   NAND2X1 U618 (.IN1(n25), .IN2(n83), .QN(n774));
   NAND2X1 U619 (.IN1(n795), .IN2(n24), .QN(n663));
   NAND2X1 U620 (.IN1(n1166), .IN2(n21), .QN(n1037));
   NAND2X1 U621 (.IN1(n18), .IN2(n241), .QN(n1303));
   NAND2X1 U622 (.IN1(n520), .IN2(n15), .QN(n422));
   NAND2X1 U623 (.IN1(n22), .IN2(n126), .QN(n1114));
   NAND2X1 U624 (.IN1(n16), .IN2(n1564), .QN(n499));
   OR2X1 U625 (.IN1(n1366), .IN2(n42), .Q(n273));
   NAND2X1 U626 (.IN1(n25), .IN2(n72), .QN(n755));
   INVX0 U627 (.INP(sboxw[23]), .ZN(n91));
   NAND2X1 U628 (.IN1(n22), .IN2(n115), .QN(n1095));
   NOR2X0 U629 (.IN1(n11), .IN2(sboxw[30]), .QN(n616));
   NAND2X1 U630 (.IN1(n16), .IN2(n1553), .QN(n480));
   NOR2X0 U631 (.IN1(n47), .IN2(sboxw[30]), .QN(n614));
   NOR2X0 U632 (.IN1(n155), .IN2(n19), .QN(n300));
   NAND2X1 U633 (.IN1(n19), .IN2(n155), .QN(n265));
   NAND2X1 U634 (.IN1(sboxw[11]), .IN2(n172), .QN(n217));
   NOR2X0 U635 (.IN1(n168), .IN2(n20), .QN(n1354));
   NAND2X1 U636 (.IN1(n1440), .IN2(n18), .QN(n1377));
   NOR2X0 U637 (.IN1(n40), .IN2(sboxw[6]), .QN(n373));
   NAND2X1 U638 (.IN1(n299), .IN2(n18), .QN(n268));
   INVX0 U639 (.INP(sboxw[3]), .ZN(n1564));
   NOR2X0 U640 (.IN1(n19), .IN2(n20), .QN(n1348));
   NAND2X1 U641 (.IN1(n25), .IN2(sboxw[27]), .QN(n638));
   INVX0 U642 (.INP(sboxw[11]), .ZN(n167));
   NOR2X0 U643 (.IN1(n48), .IN2(sboxw[30]), .QN(n545));
   INVX0 U644 (.INP(sboxw[27]), .ZN(n83));
   NAND2X1 U645 (.IN1(n16), .IN2(sboxw[3]), .QN(n397));
   NOR2X0 U646 (.IN1(n178), .IN2(sboxw[6]), .QN(n304));
   NOR2X0 U647 (.IN1(n46), .IN2(n24), .QN(n637));
   INVX0 U648 (.INP(sboxw[30]), .ZN(n49));
   NOR2X0 U649 (.IN1(n39), .IN2(n15), .QN(n396));
   NOR2X0 U650 (.IN1(n49), .IN2(n47), .QN(n550));
   INVX0 U651 (.INP(sboxw[6]), .ZN(n179));
   NOR2X0 U652 (.IN1(n9), .IN2(sboxw[14]), .QN(n1339));
   NOR2X0 U653 (.IN1(n43), .IN2(sboxw[14]), .QN(n1337));
   NOR2X0 U654 (.IN1(n134), .IN2(sboxw[14]), .QN(n1290));
   INVX0 U655 (.INP(sboxw[31]), .ZN(n48));
   INVX0 U656 (.INP(sboxw[14]), .ZN(n135));
   NOR2X0 U657 (.IN1(n135), .IN2(n9), .QN(n188));
   INVX0 U658 (.INP(n19), .ZN(n172));
   NOR2X0 U659 (.IN1(n43), .IN2(n19), .QN(n229));
   INVX0 U660 (.INP(sboxw[7]), .ZN(n178));
   INVX0 U661 (.INP(sboxw[15]), .ZN(n134));
   INVX0 U662 (.INP(n39), .ZN(n12));
   NBUFFX2 U663 (.INP(sboxw[4]), .Z(n17));
   NBUFFX2 U664 (.INP(sboxw[20]), .Z(n23));
   NBUFFX2 U665 (.INP(sboxw[28]), .Z(n26));
   INVX0 U666 (.INP(n45), .ZN(n10));
   INVX0 U667 (.INP(n40), .ZN(n8));
   INVX0 U668 (.INP(n281), .ZN(n176));
   NAND2X0 U669 (.IN1(n281), .IN2(n228), .QN(n1304));
   NOR2X0 U670 (.IN1(n179), .IN2(n8), .QN(n307));
   NOR2X0 U671 (.IN1(n8), .IN2(sboxw[6]), .QN(n375));
   NOR2X0 U672 (.IN1(n398), .IN2(n8), .QN(n440));
   OA21X1 U673 (.IN1(n331), .IN2(n1533), .IN3(n8), .Q(n1531));
   INVX0 U674 (.INP(n47), .ZN(n11));
   NOR2X0 U675 (.IN1(n47), .IN2(n25), .QN(n739));
   NAND2X0 U676 (.IN1(n708), .IN2(n47), .QN(n567));
   NAND2X0 U677 (.IN1(n87), .IN2(n47), .QN(n566));
   NOR2X0 U678 (.IN1(n172), .IN2(n9), .QN(n271));
   OA21X1 U679 (.IN1(n204), .IN2(n292), .IN3(n9), .Q(n291));
   NOR2X0 U680 (.IN1(n164), .IN2(n9), .QN(n277));
   INVX0 U681 (.INP(n43), .ZN(n9));
   INVX0 U682 (.INP(n15), .ZN(n1571));
   NOR2X0 U683 (.IN1(n33), .IN2(n572), .QN(n4));
   NOR2X0 U684 (.IN1(n33), .IN2(n572), .QN(n5));
   NOR2X0 U685 (.IN1(n35), .IN2(n331), .QN(n6));
   NOR2X0 U686 (.IN1(n35), .IN2(n331), .QN(n7));
   NOR2X0 U687 (.IN1(n39), .IN2(n181), .QN(n358));
   INVX0 U688 (.INP(n381), .ZN(n181));
   NOR2X0 U689 (.IN1(n1552), .IN2(n183), .QN(n381));
   NOR2X0 U690 (.IN1(n1547), .IN2(n183), .QN(n359));
   NOR2X0 U691 (.IN1(n1561), .IN2(n183), .QN(n317));
   INVX0 U692 (.INP(n464), .ZN(n183));
   NOR2X0 U693 (.IN1(n138), .IN2(n148), .QN(n200));
   INVX0 U694 (.INP(n996), .ZN(n94));
   NOR2X0 U695 (.IN1(n114), .IN2(n96), .QN(n996));
   NOR2X0 U696 (.IN1(n123), .IN2(n96), .QN(n932));
   NOR2X0 U697 (.IN1(n109), .IN2(n96), .QN(n974));
   INVX0 U698 (.INP(n1079), .ZN(n96));
   NOR2X0 U699 (.IN1(n45), .IN2(n22), .QN(n1079));
   NOR2X0 U700 (.IN1(n72), .IN2(sboxw[27]), .QN(n722));
   NOR2X0 U701 (.IN1(n33), .IN2(n572), .QN(n583));
   INVX0 U702 (.INP(n277), .ZN(n141));
   NOR2X0 U703 (.IN1(n172), .IN2(sboxw[11]), .QN(n299));
   NOR2X0 U704 (.IN1(n87), .IN2(n70), .QN(n813));
   INVX0 U705 (.INP(n793), .ZN(n70));
   NOR2X0 U706 (.IN1(n91), .IN2(sboxw[22]), .QN(n919));
   NOR2X0 U707 (.IN1(n45), .IN2(sboxw[22]), .QN(n988));
   NOR2X0 U708 (.IN1(n10), .IN2(sboxw[22]), .QN(n990));
   NAND2X0 U709 (.IN1(n244), .IN2(n174), .QN(n1324));
   INVX0 U710 (.INP(n1324), .ZN(n149));
   INVX0 U711 (.INP(n211), .ZN(n174));
   INVX0 U712 (.INP(sboxw[19]), .ZN(n126));
   NOR2X0 U713 (.IN1(sboxw[19]), .IN2(n23), .QN(n1006));
   NAND2X0 U714 (.IN1(sboxw[19]), .IN2(n128), .QN(n1090));
   NAND2X0 U715 (.IN1(n31), .IN2(sboxw[19]), .QN(n1031));
   OA21X1 U716 (.IN1(n23), .IN2(n1011), .IN3(sboxw[19]), .Q(n1030));
   NOR2X0 U717 (.IN1(n1001), .IN2(n1002), .QN(n999));
   NOR2X0 U718 (.IN1(n128), .IN2(n109), .QN(n1002));
   NOR2X0 U719 (.IN1(n115), .IN2(sboxw[19]), .QN(n1062));
   NOR2X0 U720 (.IN1(n1013), .IN2(n10), .QN(n1055));
   INVX0 U721 (.INP(n1164), .ZN(n113));
   NAND2X0 U722 (.IN1(n1164), .IN2(n21), .QN(n1024));
   INVX0 U723 (.INP(n937), .ZN(n117));
   NOR2X0 U724 (.IN1(n128), .IN2(n114), .QN(n1164));
   INVX0 U725 (.INP(n2), .ZN(n34));
   INVX0 U726 (.INP(n44), .ZN(n13));
   NOR2X0 U727 (.IN1(n35), .IN2(n331), .QN(n342));
   OA21X1 U728 (.IN1(n148), .IN2(n41), .IN3(n147), .Q(n234));
   NAND2X0 U729 (.IN1(n245), .IN2(n42), .QN(n1351));
   OA21X1 U730 (.IN1(n41), .IN2(n162), .IN3(n213), .Q(n1373));
   NAND2X0 U731 (.IN1(n1355), .IN2(n41), .QN(n1442));
   NAND2X0 U732 (.IN1(n41), .IN2(n1349), .QN(n207));
   NAND2X0 U733 (.IN1(n206), .IN2(n42), .QN(n1505));
   NAND2X0 U734 (.IN1(n228), .IN2(n41), .QN(n1311));
   NAND2X0 U735 (.IN1(n200), .IN2(n41), .QN(n1318));
   NAND2X0 U736 (.IN1(n41), .IN2(n250), .QN(n1302));
   NAND2X0 U737 (.IN1(n242), .IN2(n42), .QN(n1325));
   NAND2X0 U738 (.IN1(n1375), .IN2(n41), .QN(n225));
   NOR2X0 U739 (.IN1(n152), .IN2(n42), .QN(n262));
   NOR2X0 U740 (.IN1(n41), .IN2(n18), .QN(n204));
   NOR2X0 U741 (.IN1(n42), .IN2(n18), .QN(n201));
   NOR2X0 U742 (.IN1(n177), .IN2(n41), .QN(n281));
   INVX0 U743 (.INP(n32), .ZN(n31));
   INVX0 U744 (.INP(n46), .ZN(n14));
   NOR2X0 U745 (.IN1(n19), .IN2(n9), .QN(n286));
   INVX0 U746 (.INP(n3), .ZN(n38));
   INVX0 U747 (.INP(n3), .ZN(n37));
   INVX0 U748 (.INP(n24), .ZN(n90));
   INVX0 U749 (.INP(sboxw[21]), .ZN(n45));
   INVX0 U750 (.INP(sboxw[1]), .ZN(n39));
   NOR2X0 U751 (.IN1(n356), .IN2(n518), .QN(n528));
   NOR2X0 U752 (.IN1(n446), .IN2(n356), .QN(n463));
   INVX0 U826 (.INP(sboxw[5]), .ZN(n40));
   NAND2X0 U829 (.IN1(n360), .IN2(n361), .QN(n303));
   NOR2X0 U853 (.IN1(n1540), .IN2(n1564), .QN(n684));
   INVX0 U890 (.INP(n405), .ZN(n185));
   NOR2X0 U903 (.IN1(n205), .IN2(n396), .QN(n405));
   NOR2X0 U931 (.IN1(n1557), .IN2(n323), .QN(n460));
   INVX0 U956 (.INP(n460), .ZN(n184));
   INVX0 U980 (.INP(sboxw[25]), .ZN(n46));
   OA21X1 U994 (.IN1(n1570), .IN2(n205), .IN3(n363), .Q(n533));
   INVX0 U1025 (.INP(n327), .ZN(n1540));
   NOR2X0 U1104 (.IN1(n40), .IN2(n16), .QN(n464));
   NOR2X0 U1165 (.IN1(n323), .IN2(n1552), .QN(n542));
   NAND2X0 U1167 (.IN1(n542), .IN2(n35), .QN(n363));
   INVX0 U1172 (.INP(sboxw[9]), .ZN(n42));
   INVX0 U1188 (.INP(n1519), .ZN(n205));
   NOR2X0 U1208 (.IN1(n323), .IN2(n1547), .QN(n1519));
   INVX0 U1214 (.INP(n286), .ZN(n143));
   INVX0 U1215 (.INP(sboxw[13]), .ZN(n43));
   NAND2X0 U1233 (.IN1(n269), .IN2(n37), .QN(n1329));
   NAND2X0 U1242 (.IN1(n269), .IN2(n211), .QN(n274));
   NAND2X1 U1244 (.IN1(n269), .IN2(n18), .QN(n256));
   NOR2X0 U1245 (.IN1(n143), .IN2(n148), .QN(n269));
   NOR2X0 U1258 (.IN1(n76), .IN2(n57), .QN(n735));
   INVX0 U1289 (.INP(sboxw[29]), .ZN(n47));
   INVX0 U1317 (.INP(n1), .ZN(n36));
   NAND2X0 U1333 (.IN1(n131), .IN2(n1016), .QN(n1025));
   INVX0 U1352 (.INP(sboxw[17]), .ZN(n44));
   INVX0 U1368 (.INP(n946), .ZN(n131));
   NOR2X0 U1381 (.IN1(n133), .IN2(n13), .QN(n985));
   OA21X1 U1386 (.IN1(n946), .IN2(n108), .IN3(n1008), .Q(n1285));
   OA21X1 U1393 (.IN1(n946), .IN2(n1281), .IN3(n10), .Q(n1279));
   NAND2X0 U1396 (.IN1(n946), .IN2(n1006), .QN(n961));
   NAND2X0 U1427 (.IN1(n1006), .IN2(n957), .QN(n1049));
   NAND2X0 U1514 (.IN1(n946), .IN2(n128), .QN(n1007));
   NAND2X0 U1519 (.IN1(n937), .IN2(n957), .QN(n1038));
   NAND2X0 U1521 (.IN1(n1164), .IN2(n957), .QN(n1057));
   OA21X1 U1536 (.IN1(n117), .IN2(n946), .IN3(n936), .Q(n983));
   NOR2X0 U1542 (.IN1(n947), .IN2(n132), .QN(n1047));
   INVX0 U1546 (.INP(n985), .ZN(n132));
   OA21X1 U1549 (.IN1(sboxw[17]), .IN2(n120), .IN3(n969), .Q(n1033));
   NOR2X0 U1556 (.IN1(n938), .IN2(n946), .QN(n957));
   NOR2X0 U1572 (.IN1(n13), .IN2(n21), .QN(n946));
   NOR2X0 U1573 (.IN1(n128), .IN2(n10), .QN(n942));
   NAND2X0 U1574 (.IN1(n518), .IN2(n1567), .QN(n354));
   NAND2X0 U1575 (.IN1(n541), .IN2(n1567), .QN(n393));
   NAND2X0 U1576 (.IN1(n387), .IN2(n1567), .QN(n454));
   NOR2X0 U1577 (.IN1(n1567), .IN2(n1552), .QN(n356));
   INVX0 U1578 (.INP(n957), .ZN(n129));
   NOR2X0 U1579 (.IN1(n1566), .IN2(n8), .QN(n327));
   INVX0 U1580 (.INP(n366), .ZN(n323));
   NOR2X0 U1581 (.IN1(n16), .IN2(n8), .QN(n366));
   INVX0 U1582 (.INP(n981), .ZN(n100));
   NOR2X0 U1583 (.IN1(n22), .IN2(n10), .QN(n981));
   NAND2X0 U1584 (.IN1(n793), .IN2(n86), .QN(n595));
   NAND2X0 U1585 (.IN1(n816), .IN2(n86), .QN(n634));
   NAND2X0 U1586 (.IN1(n628), .IN2(n86), .QN(n729));
   NOR2X0 U1587 (.IN1(n86), .IN2(n71), .QN(n597));
   NOR2X0 U1588 (.IN1(n971), .IN2(n1164), .QN(n1174));
   NOR2X0 U1589 (.IN1(n1061), .IN2(n971), .QN(n1078));
   NOR2X0 U1590 (.IN1(n133), .IN2(n44), .QN(n938));
   NAND2X0 U1591 (.IN1(n1188), .IN2(n129), .QN(n1269));
   NAND2X0 U1592 (.IN1(n931), .IN2(n129), .QN(n1161));
   OA21X1 U1593 (.IN1(n129), .IN2(n120), .IN3(n983), .Q(n1215));
   NAND2X0 U1594 (.IN1(n1048), .IN2(n129), .QN(n1243));
   OA21X1 U1595 (.IN1(n931), .IN2(n937), .IN3(n129), .Q(n1178));
   NOR2X0 U1596 (.IN1(n129), .IN2(n114), .QN(n971));
   NAND2X0 U1597 (.IN1(n1002), .IN2(n129), .QN(n1069));
   NAND2X0 U1598 (.IN1(n1187), .IN2(n129), .QN(n1008));
   NAND2X0 U1599 (.IN1(n1164), .IN2(n129), .QN(n969));
   NBUFFX2 U1600 (.INP(n201), .Z(n27));
   NBUFFX2 U1601 (.INP(n201), .Z(n28));
   NBUFFX2 U1602 (.INP(n201), .Z(n29));
   NBUFFX2 U1603 (.INP(n201), .Z(n30));
endmodule

module aes_core_test_1 (clk, reset_n, encdec, init, next, ready, key, keylen, block, 
       result, result_valid, test_si3, test_si2, test_si1, test_so3, test_so2, test_so1, 
       test_se);
input clk, reset_n, encdec, init, next, keylen, test_si3, test_si2, test_si1, test_se;
input [255:0] key;
input [127:0] block;
output ready, result_valid, test_so3, test_so2, test_so1;
output [127:0] result;
wire enc_next, enc_ready, dec_next, dec_ready, key_ready, n6, n9, n12, n13, n14, n15, n16
       , n17, n18, n19, n20, n21, n23, n24, n25, n26, n5, n7, n8, n10, n11, n22, n27, n28
       , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, 
       n45, n46, n47, n48, n49, n52, n53, n56, n57;
wire [3:0] enc_round_nr;
wire [127:0] round_key;
wire [31:0] enc_sboxw;
wire [31:0] new_sboxw;
wire [127:0] enc_new_block;
wire [3:0] dec_round_nr;
wire [127:0] dec_new_block;
wire [3:0] muxed_round_nr;
wire [31:0] keymem_sboxw;
wire [31:0] muxed_sboxw;
wire [1:0] aes_core_ctrl_reg;
   SDFFARX1 \aes_core_ctrl_reg_reg[0]  (.D(n26), .SI(test_si1), .SE(test_se), .CLK(clk), .
          RSTB(n45), .Q(aes_core_ctrl_reg[0]), .QN(n9));
   SDFFASX1 ready_reg_reg (.D(n24), .SI(n53), .SE(test_se), .CLK(clk), .SETB(n45), .Q(
          ready), .QN(n52));
   SDFFARX1 result_valid_reg_reg (.D(n23), .SI(n52), .SE(test_se), .CLK(clk), .RSTB(n45), .
          Q(result_valid), .QN(test_so3));
   AO22X1 U20 (.IN1(n11), .IN2(enc_new_block[9]), .IN3(dec_new_block[9]), .IN4(n36), .Q(
          result[9]));
   AO22X1 U21 (.IN1(enc_new_block[99]), .IN2(n11), .IN3(dec_new_block[99]), .IN4(n36), .Q(
          result[99]));
   AO22X1 U22 (.IN1(enc_new_block[98]), .IN2(n11), .IN3(dec_new_block[98]), .IN4(n36), .Q(
          result[98]));
   AO22X1 U23 (.IN1(enc_new_block[97]), .IN2(n11), .IN3(dec_new_block[97]), .IN4(n36), .Q(
          result[97]));
   AO22X1 U24 (.IN1(enc_new_block[96]), .IN2(n11), .IN3(dec_new_block[96]), .IN4(n36), .Q(
          result[96]));
   AO22X1 U25 (.IN1(enc_new_block[95]), .IN2(n11), .IN3(dec_new_block[95]), .IN4(n36), .Q(
          result[95]));
   AO22X1 U26 (.IN1(enc_new_block[94]), .IN2(n11), .IN3(dec_new_block[94]), .IN4(n36), .Q(
          result[94]));
   AO22X1 U27 (.IN1(enc_new_block[93]), .IN2(n11), .IN3(dec_new_block[93]), .IN4(n36), .Q(
          result[93]));
   AO22X1 U28 (.IN1(enc_new_block[92]), .IN2(n11), .IN3(dec_new_block[92]), .IN4(n36), .Q(
          result[92]));
   AO22X1 U29 (.IN1(enc_new_block[91]), .IN2(n11), .IN3(dec_new_block[91]), .IN4(n36), .Q(
          result[91]));
   AO22X1 U30 (.IN1(enc_new_block[90]), .IN2(n11), .IN3(dec_new_block[90]), .IN4(n36), .Q(
          result[90]));
   AO22X1 U31 (.IN1(enc_new_block[8]), .IN2(n11), .IN3(dec_new_block[8]), .IN4(n36), .Q(
          result[8]));
   AO22X1 U32 (.IN1(enc_new_block[89]), .IN2(n11), .IN3(dec_new_block[89]), .IN4(n36), .Q(
          result[89]));
   AO22X1 U33 (.IN1(enc_new_block[88]), .IN2(n11), .IN3(dec_new_block[88]), .IN4(n36), .Q(
          result[88]));
   AO22X1 U34 (.IN1(enc_new_block[87]), .IN2(n11), .IN3(dec_new_block[87]), .IN4(n36), .Q(
          result[87]));
   AO22X1 U35 (.IN1(enc_new_block[86]), .IN2(n22), .IN3(dec_new_block[86]), .IN4(n36), .Q(
          result[86]));
   AO22X1 U36 (.IN1(enc_new_block[85]), .IN2(n22), .IN3(dec_new_block[85]), .IN4(n36), .Q(
          result[85]));
   AO22X1 U37 (.IN1(enc_new_block[84]), .IN2(n22), .IN3(dec_new_block[84]), .IN4(n36), .Q(
          result[84]));
   AO22X1 U38 (.IN1(enc_new_block[83]), .IN2(n22), .IN3(dec_new_block[83]), .IN4(n36), .Q(
          result[83]));
   AO22X1 U39 (.IN1(enc_new_block[82]), .IN2(n22), .IN3(dec_new_block[82]), .IN4(n36), .Q(
          result[82]));
   AO22X1 U40 (.IN1(enc_new_block[81]), .IN2(n22), .IN3(dec_new_block[81]), .IN4(n36), .Q(
          result[81]));
   AO22X1 U41 (.IN1(enc_new_block[80]), .IN2(n22), .IN3(dec_new_block[80]), .IN4(n36), .Q(
          result[80]));
   AO22X1 U42 (.IN1(enc_new_block[7]), .IN2(n22), .IN3(dec_new_block[7]), .IN4(n36), .Q(
          result[7]));
   AO22X1 U43 (.IN1(enc_new_block[79]), .IN2(n22), .IN3(dec_new_block[79]), .IN4(n36), .Q(
          result[79]));
   AO22X1 U44 (.IN1(enc_new_block[78]), .IN2(n22), .IN3(dec_new_block[78]), .IN4(n36), .Q(
          result[78]));
   AO22X1 U45 (.IN1(enc_new_block[77]), .IN2(n22), .IN3(dec_new_block[77]), .IN4(n36), .Q(
          result[77]));
   AO22X1 U46 (.IN1(enc_new_block[76]), .IN2(n22), .IN3(dec_new_block[76]), .IN4(n36), .Q(
          result[76]));
   AO22X1 U47 (.IN1(enc_new_block[75]), .IN2(n22), .IN3(dec_new_block[75]), .IN4(n36), .Q(
          result[75]));
   AO22X1 U48 (.IN1(enc_new_block[74]), .IN2(n22), .IN3(dec_new_block[74]), .IN4(n36), .Q(
          result[74]));
   AO22X1 U49 (.IN1(enc_new_block[73]), .IN2(n22), .IN3(dec_new_block[73]), .IN4(n36), .Q(
          result[73]));
   AO22X1 U50 (.IN1(enc_new_block[72]), .IN2(n22), .IN3(dec_new_block[72]), .IN4(n36), .Q(
          result[72]));
   AO22X1 U51 (.IN1(enc_new_block[71]), .IN2(n22), .IN3(dec_new_block[71]), .IN4(n36), .Q(
          result[71]));
   AO22X1 U52 (.IN1(enc_new_block[70]), .IN2(n27), .IN3(dec_new_block[70]), .IN4(n37), .Q(
          result[70]));
   AO22X1 U53 (.IN1(enc_new_block[6]), .IN2(n27), .IN3(dec_new_block[6]), .IN4(n37), .Q(
          result[6]));
   AO22X1 U54 (.IN1(enc_new_block[69]), .IN2(n27), .IN3(dec_new_block[69]), .IN4(n37), .Q(
          result[69]));
   AO22X1 U55 (.IN1(enc_new_block[68]), .IN2(n27), .IN3(dec_new_block[68]), .IN4(n37), .Q(
          result[68]));
   AO22X1 U56 (.IN1(enc_new_block[67]), .IN2(n27), .IN3(dec_new_block[67]), .IN4(n37), .Q(
          result[67]));
   AO22X1 U57 (.IN1(enc_new_block[66]), .IN2(n27), .IN3(dec_new_block[66]), .IN4(n37), .Q(
          result[66]));
   AO22X1 U58 (.IN1(enc_new_block[65]), .IN2(n27), .IN3(dec_new_block[65]), .IN4(n37), .Q(
          result[65]));
   AO22X1 U59 (.IN1(enc_new_block[64]), .IN2(n27), .IN3(dec_new_block[64]), .IN4(n37), .Q(
          result[64]));
   AO22X1 U60 (.IN1(enc_new_block[63]), .IN2(n27), .IN3(dec_new_block[63]), .IN4(n37), .Q(
          result[63]));
   AO22X1 U61 (.IN1(enc_new_block[62]), .IN2(n27), .IN3(dec_new_block[62]), .IN4(n37), .Q(
          result[62]));
   AO22X1 U62 (.IN1(enc_new_block[61]), .IN2(n27), .IN3(dec_new_block[61]), .IN4(n37), .Q(
          result[61]));
   AO22X1 U63 (.IN1(enc_new_block[60]), .IN2(n27), .IN3(dec_new_block[60]), .IN4(n37), .Q(
          result[60]));
   AO22X1 U64 (.IN1(enc_new_block[5]), .IN2(n27), .IN3(dec_new_block[5]), .IN4(n38), .Q(
          result[5]));
   AO22X1 U65 (.IN1(enc_new_block[59]), .IN2(n27), .IN3(dec_new_block[59]), .IN4(n38), .Q(
          result[59]));
   AO22X1 U66 (.IN1(enc_new_block[58]), .IN2(n27), .IN3(dec_new_block[58]), .IN4(n38), .Q(
          result[58]));
   AO22X1 U67 (.IN1(enc_new_block[57]), .IN2(n27), .IN3(dec_new_block[57]), .IN4(n38), .Q(
          result[57]));
   AO22X1 U68 (.IN1(enc_new_block[56]), .IN2(n27), .IN3(dec_new_block[56]), .IN4(n38), .Q(
          result[56]));
   AO22X1 U69 (.IN1(enc_new_block[55]), .IN2(n28), .IN3(dec_new_block[55]), .IN4(n38), .Q(
          result[55]));
   AO22X1 U70 (.IN1(enc_new_block[54]), .IN2(n28), .IN3(dec_new_block[54]), .IN4(n38), .Q(
          result[54]));
   AO22X1 U71 (.IN1(enc_new_block[53]), .IN2(n28), .IN3(dec_new_block[53]), .IN4(n38), .Q(
          result[53]));
   AO22X1 U72 (.IN1(enc_new_block[52]), .IN2(n28), .IN3(dec_new_block[52]), .IN4(n38), .Q(
          result[52]));
   AO22X1 U73 (.IN1(enc_new_block[51]), .IN2(n28), .IN3(dec_new_block[51]), .IN4(n38), .Q(
          result[51]));
   AO22X1 U74 (.IN1(enc_new_block[50]), .IN2(n28), .IN3(dec_new_block[50]), .IN4(n38), .Q(
          result[50]));
   AO22X1 U75 (.IN1(enc_new_block[4]), .IN2(n28), .IN3(dec_new_block[4]), .IN4(n38), .Q(
          result[4]));
   AO22X1 U76 (.IN1(enc_new_block[49]), .IN2(n28), .IN3(dec_new_block[49]), .IN4(n39), .Q(
          result[49]));
   AO22X1 U77 (.IN1(enc_new_block[48]), .IN2(n28), .IN3(dec_new_block[48]), .IN4(n39), .Q(
          result[48]));
   AO22X1 U78 (.IN1(enc_new_block[47]), .IN2(n28), .IN3(dec_new_block[47]), .IN4(n39), .Q(
          result[47]));
   AO22X1 U79 (.IN1(enc_new_block[46]), .IN2(n28), .IN3(dec_new_block[46]), .IN4(n39), .Q(
          result[46]));
   AO22X1 U80 (.IN1(enc_new_block[45]), .IN2(n28), .IN3(dec_new_block[45]), .IN4(n39), .Q(
          result[45]));
   AO22X1 U81 (.IN1(enc_new_block[44]), .IN2(n28), .IN3(dec_new_block[44]), .IN4(n39), .Q(
          result[44]));
   AO22X1 U82 (.IN1(enc_new_block[43]), .IN2(n28), .IN3(dec_new_block[43]), .IN4(n39), .Q(
          result[43]));
   AO22X1 U83 (.IN1(enc_new_block[42]), .IN2(n28), .IN3(dec_new_block[42]), .IN4(n39), .Q(
          result[42]));
   AO22X1 U84 (.IN1(enc_new_block[41]), .IN2(n28), .IN3(dec_new_block[41]), .IN4(n39), .Q(
          result[41]));
   AO22X1 U85 (.IN1(enc_new_block[40]), .IN2(n28), .IN3(dec_new_block[40]), .IN4(n39), .Q(
          result[40]));
   AO22X1 U86 (.IN1(enc_new_block[3]), .IN2(n29), .IN3(dec_new_block[3]), .IN4(n39), .Q(
          result[3]));
   AO22X1 U87 (.IN1(enc_new_block[39]), .IN2(n29), .IN3(dec_new_block[39]), .IN4(n44), .Q(
          result[39]));
   AO22X1 U88 (.IN1(enc_new_block[38]), .IN2(n29), .IN3(dec_new_block[38]), .IN4(n44), .Q(
          result[38]));
   AO22X1 U89 (.IN1(enc_new_block[37]), .IN2(n29), .IN3(dec_new_block[37]), .IN4(n44), .Q(
          result[37]));
   AO22X1 U90 (.IN1(enc_new_block[36]), .IN2(n29), .IN3(dec_new_block[36]), .IN4(n44), .Q(
          result[36]));
   AO22X1 U91 (.IN1(enc_new_block[35]), .IN2(n29), .IN3(dec_new_block[35]), .IN4(n44), .Q(
          result[35]));
   AO22X1 U92 (.IN1(enc_new_block[34]), .IN2(n29), .IN3(dec_new_block[34]), .IN4(n44), .Q(
          result[34]));
   AO22X1 U93 (.IN1(enc_new_block[33]), .IN2(n29), .IN3(dec_new_block[33]), .IN4(n44), .Q(
          result[33]));
   AO22X1 U94 (.IN1(enc_new_block[32]), .IN2(n29), .IN3(dec_new_block[32]), .IN4(n44), .Q(
          result[32]));
   AO22X1 U95 (.IN1(enc_new_block[31]), .IN2(n29), .IN3(dec_new_block[31]), .IN4(n44), .Q(
          result[31]));
   AO22X1 U96 (.IN1(enc_new_block[30]), .IN2(n29), .IN3(dec_new_block[30]), .IN4(n44), .Q(
          result[30]));
   AO22X1 U97 (.IN1(enc_new_block[2]), .IN2(n29), .IN3(dec_new_block[2]), .IN4(n44), .Q(
          result[2]));
   AO22X1 U98 (.IN1(enc_new_block[29]), .IN2(n29), .IN3(dec_new_block[29]), .IN4(n44), .Q(
          result[29]));
   AO22X1 U99 (.IN1(enc_new_block[28]), .IN2(n29), .IN3(dec_new_block[28]), .IN4(n44), .Q(
          result[28]));
   AO22X1 U100 (.IN1(enc_new_block[27]), .IN2(n29), .IN3(dec_new_block[27]), .IN4(n44), .Q(
          result[27]));
   AO22X1 U101 (.IN1(enc_new_block[26]), .IN2(n29), .IN3(dec_new_block[26]), .IN4(n44), .Q(
          result[26]));
   AO22X1 U102 (.IN1(enc_new_block[25]), .IN2(n29), .IN3(dec_new_block[25]), .IN4(n44), .Q(
          result[25]));
   AO22X1 U103 (.IN1(enc_new_block[24]), .IN2(n30), .IN3(dec_new_block[24]), .IN4(n44), .Q(
          result[24]));
   AO22X1 U104 (.IN1(enc_new_block[23]), .IN2(n30), .IN3(dec_new_block[23]), .IN4(n44), .Q(
          result[23]));
   AO22X1 U105 (.IN1(enc_new_block[22]), .IN2(n30), .IN3(dec_new_block[22]), .IN4(n44), .Q(
          result[22]));
   AO22X1 U106 (.IN1(enc_new_block[21]), .IN2(n30), .IN3(dec_new_block[21]), .IN4(n44), .Q(
          result[21]));
   AO22X1 U107 (.IN1(enc_new_block[20]), .IN2(n30), .IN3(dec_new_block[20]), .IN4(n44), .Q(
          result[20]));
   AO22X1 U108 (.IN1(enc_new_block[1]), .IN2(n30), .IN3(dec_new_block[1]), .IN4(n44), .Q(
          result[1]));
   AO22X1 U109 (.IN1(enc_new_block[19]), .IN2(n30), .IN3(dec_new_block[19]), .IN4(n40), .Q(
          result[19]));
   AO22X1 U110 (.IN1(enc_new_block[18]), .IN2(n30), .IN3(dec_new_block[18]), .IN4(n40), .Q(
          result[18]));
   AO22X1 U111 (.IN1(enc_new_block[17]), .IN2(n30), .IN3(dec_new_block[17]), .IN4(n40), .Q(
          result[17]));
   AO22X1 U112 (.IN1(enc_new_block[16]), .IN2(n30), .IN3(dec_new_block[16]), .IN4(n40), .Q(
          result[16]));
   AO22X1 U113 (.IN1(enc_new_block[15]), .IN2(n30), .IN3(dec_new_block[15]), .IN4(n40), .Q(
          result[15]));
   AO22X1 U114 (.IN1(enc_new_block[14]), .IN2(n30), .IN3(dec_new_block[14]), .IN4(n40), .Q(
          result[14]));
   AO22X1 U115 (.IN1(enc_new_block[13]), .IN2(n30), .IN3(dec_new_block[13]), .IN4(n40), .Q(
          result[13]));
   AO22X1 U116 (.IN1(enc_new_block[12]), .IN2(n30), .IN3(dec_new_block[12]), .IN4(n40), .Q(
          result[12]));
   AO22X1 U117 (.IN1(enc_new_block[127]), .IN2(n30), .IN3(dec_new_block[127]), .IN4(n40), .
          Q(result[127]));
   AO22X1 U118 (.IN1(enc_new_block[126]), .IN2(n30), .IN3(dec_new_block[126]), .IN4(n40), .
          Q(result[126]));
   AO22X1 U119 (.IN1(enc_new_block[125]), .IN2(n30), .IN3(dec_new_block[125]), .IN4(n40), .
          Q(result[125]));
   AO22X1 U120 (.IN1(enc_new_block[124]), .IN2(n31), .IN3(dec_new_block[124]), .IN4(n40), .
          Q(result[124]));
   AO22X1 U121 (.IN1(enc_new_block[123]), .IN2(n31), .IN3(dec_new_block[123]), .IN4(n39), .
          Q(result[123]));
   AO22X1 U122 (.IN1(enc_new_block[122]), .IN2(n31), .IN3(dec_new_block[122]), .IN4(n41), .
          Q(result[122]));
   AO22X1 U123 (.IN1(enc_new_block[121]), .IN2(n31), .IN3(dec_new_block[121]), .IN4(n41), .
          Q(result[121]));
   AO22X1 U124 (.IN1(enc_new_block[120]), .IN2(n31), .IN3(dec_new_block[120]), .IN4(n41), .
          Q(result[120]));
   AO22X1 U125 (.IN1(enc_new_block[11]), .IN2(n31), .IN3(dec_new_block[11]), .IN4(n41), .Q(
          result[11]));
   AO22X1 U126 (.IN1(enc_new_block[119]), .IN2(n31), .IN3(dec_new_block[119]), .IN4(n41), .
          Q(result[119]));
   AO22X1 U127 (.IN1(enc_new_block[118]), .IN2(n31), .IN3(dec_new_block[118]), .IN4(n41), .
          Q(result[118]));
   AO22X1 U128 (.IN1(enc_new_block[117]), .IN2(n31), .IN3(dec_new_block[117]), .IN4(n41), .
          Q(result[117]));
   AO22X1 U129 (.IN1(enc_new_block[116]), .IN2(n31), .IN3(dec_new_block[116]), .IN4(n41), .
          Q(result[116]));
   AO22X1 U130 (.IN1(enc_new_block[115]), .IN2(n31), .IN3(dec_new_block[115]), .IN4(n41), .
          Q(result[115]));
   AO22X1 U131 (.IN1(enc_new_block[114]), .IN2(n31), .IN3(dec_new_block[114]), .IN4(n41), .
          Q(result[114]));
   AO22X1 U132 (.IN1(enc_new_block[113]), .IN2(n31), .IN3(dec_new_block[113]), .IN4(n41), .
          Q(result[113]));
   AO22X1 U133 (.IN1(enc_new_block[112]), .IN2(n31), .IN3(dec_new_block[112]), .IN4(n41), .
          Q(result[112]));
   AO22X1 U134 (.IN1(enc_new_block[111]), .IN2(n31), .IN3(dec_new_block[111]), .IN4(n43), .
          Q(result[111]));
   AO22X1 U135 (.IN1(enc_new_block[110]), .IN2(n31), .IN3(dec_new_block[110]), .IN4(n43), .
          Q(result[110]));
   AO22X1 U136 (.IN1(enc_new_block[10]), .IN2(n31), .IN3(dec_new_block[10]), .IN4(n43), .Q(
          result[10]));
   AO22X1 U137 (.IN1(enc_new_block[109]), .IN2(n32), .IN3(dec_new_block[109]), .IN4(n41), .
          Q(result[109]));
   AO22X1 U138 (.IN1(enc_new_block[108]), .IN2(n32), .IN3(dec_new_block[108]), .IN4(n43), .
          Q(result[108]));
   AO22X1 U139 (.IN1(enc_new_block[107]), .IN2(n32), .IN3(dec_new_block[107]), .IN4(n43), .
          Q(result[107]));
   AO22X1 U140 (.IN1(enc_new_block[106]), .IN2(n32), .IN3(dec_new_block[106]), .IN4(n43), .
          Q(result[106]));
   AO22X1 U141 (.IN1(enc_new_block[105]), .IN2(n32), .IN3(dec_new_block[105]), .IN4(n43), .
          Q(result[105]));
   AO22X1 U142 (.IN1(enc_new_block[104]), .IN2(n32), .IN3(dec_new_block[104]), .IN4(n43), .
          Q(result[104]));
   AO22X1 U143 (.IN1(enc_new_block[103]), .IN2(n32), .IN3(dec_new_block[103]), .IN4(n43), .
          Q(result[103]));
   AO22X1 U144 (.IN1(enc_new_block[102]), .IN2(encdec), .IN3(dec_new_block[102]), .IN4(n43)
          , .Q(result[102]));
   AO22X1 U145 (.IN1(enc_new_block[101]), .IN2(encdec), .IN3(dec_new_block[101]), .IN4(n41)
          , .Q(result[101]));
   AO22X1 U146 (.IN1(enc_new_block[100]), .IN2(encdec), .IN3(dec_new_block[100]), .IN4(n39)
          , .Q(result[100]));
   AO22X1 U147 (.IN1(enc_new_block[0]), .IN2(encdec), .IN3(dec_new_block[0]), .IN4(n38), .
          Q(result[0]));
   AO21X1 U148 (.IN1(result_valid), .IN2(n12), .IN3(n47), .Q(n23));
   NAND3X0 U149 (.IN1(n13), .IN2(n14), .IN3(n15), .QN(n24));
   AO21X1 U151 (.IN1(n16), .IN2(aes_core_ctrl_reg[0]), .IN3(n48), .Q(n26));
   AND2X1 U152 (.IN1(n12), .IN2(n14), .Q(n16));
   NAND3X0 U153 (.IN1(aes_core_ctrl_reg[0]), .IN2(n6), .IN3(key_ready), .QN(n14));
   AO22X1 U156 (.IN1(enc_ready), .IN2(encdec), .IN3(dec_ready), .IN4(n37), .Q(n21));
   AO22X1 U157 (.IN1(keymem_sboxw[9]), .IN2(n10), .IN3(enc_sboxw[9]), .IN4(n7), .Q(
          muxed_sboxw[9]));
   AO22X1 U158 (.IN1(keymem_sboxw[8]), .IN2(n42), .IN3(enc_sboxw[8]), .IN4(n5), .Q(
          muxed_sboxw[8]));
   AO22X1 U159 (.IN1(keymem_sboxw[7]), .IN2(n10), .IN3(enc_sboxw[7]), .IN4(n5), .Q(
          muxed_sboxw[7]));
   AO22X1 U160 (.IN1(keymem_sboxw[6]), .IN2(n10), .IN3(enc_sboxw[6]), .IN4(n7), .Q(
          muxed_sboxw[6]));
   AO22X1 U162 (.IN1(keymem_sboxw[4]), .IN2(n42), .IN3(enc_sboxw[4]), .IN4(n5), .Q(
          muxed_sboxw[4]));
   AO22X1 U163 (.IN1(keymem_sboxw[3]), .IN2(n10), .IN3(enc_sboxw[3]), .IN4(n7), .Q(
          muxed_sboxw[3]));
   AO22X1 U164 (.IN1(keymem_sboxw[31]), .IN2(n42), .IN3(enc_sboxw[31]), .IN4(n7), .Q(
          muxed_sboxw[31]));
   AO22X1 U165 (.IN1(keymem_sboxw[30]), .IN2(n10), .IN3(enc_sboxw[30]), .IN4(n7), .Q(
          muxed_sboxw[30]));
   AO22X1 U166 (.IN1(keymem_sboxw[2]), .IN2(n42), .IN3(enc_sboxw[2]), .IN4(n5), .Q(
          muxed_sboxw[2]));
   AO22X1 U168 (.IN1(keymem_sboxw[28]), .IN2(n42), .IN3(enc_sboxw[28]), .IN4(n5), .Q(
          muxed_sboxw[28]));
   AO22X1 U169 (.IN1(keymem_sboxw[27]), .IN2(n42), .IN3(enc_sboxw[27]), .IN4(n7), .Q(
          muxed_sboxw[27]));
   AO22X1 U170 (.IN1(keymem_sboxw[26]), .IN2(n42), .IN3(enc_sboxw[26]), .IN4(n5), .Q(
          muxed_sboxw[26]));
   AO22X1 U171 (.IN1(keymem_sboxw[25]), .IN2(n42), .IN3(enc_sboxw[25]), .IN4(n7), .Q(
          muxed_sboxw[25]));
   AO22X1 U172 (.IN1(keymem_sboxw[24]), .IN2(n42), .IN3(enc_sboxw[24]), .IN4(n5), .Q(
          muxed_sboxw[24]));
   AO22X1 U173 (.IN1(keymem_sboxw[23]), .IN2(n42), .IN3(enc_sboxw[23]), .IN4(n7), .Q(
          muxed_sboxw[23]));
   AO22X1 U175 (.IN1(keymem_sboxw[21]), .IN2(n10), .IN3(enc_sboxw[21]), .IN4(n7), .Q(
          muxed_sboxw[21]));
   AO22X1 U176 (.IN1(keymem_sboxw[20]), .IN2(n10), .IN3(enc_sboxw[20]), .IN4(n7), .Q(
          muxed_sboxw[20]));
   AO22X1 U177 (.IN1(keymem_sboxw[1]), .IN2(n42), .IN3(enc_sboxw[1]), .IN4(n7), .Q(
          muxed_sboxw[1]));
   AO22X1 U179 (.IN1(keymem_sboxw[18]), .IN2(n10), .IN3(enc_sboxw[18]), .IN4(n7), .Q(
          muxed_sboxw[18]));
   AO22X1 U181 (.IN1(keymem_sboxw[16]), .IN2(n42), .IN3(enc_sboxw[16]), .IN4(n5), .Q(
          muxed_sboxw[16]));
   AO22X1 U182 (.IN1(keymem_sboxw[15]), .IN2(n10), .IN3(enc_sboxw[15]), .IN4(n5), .Q(
          muxed_sboxw[15]));
   AO22X1 U183 (.IN1(keymem_sboxw[14]), .IN2(n10), .IN3(enc_sboxw[14]), .IN4(n5), .Q(
          muxed_sboxw[14]));
   AO22X1 U185 (.IN1(keymem_sboxw[12]), .IN2(n42), .IN3(enc_sboxw[12]), .IN4(n5), .Q(
          muxed_sboxw[12]));
   AO22X1 U186 (.IN1(keymem_sboxw[11]), .IN2(n10), .IN3(enc_sboxw[11]), .IN4(n7), .Q(
          muxed_sboxw[11]));
   AO22X1 U187 (.IN1(keymem_sboxw[10]), .IN2(n10), .IN3(enc_sboxw[10]), .IN4(n5), .Q(
          muxed_sboxw[10]));
   AO22X1 U188 (.IN1(keymem_sboxw[0]), .IN2(n42), .IN3(enc_sboxw[0]), .IN4(n5), .Q(
          muxed_sboxw[0]));
   AO22X1 U189 (.IN1(enc_round_nr[3]), .IN2(encdec), .IN3(dec_round_nr[3]), .IN4(n43), .Q(
          muxed_round_nr[3]));
   AO22X1 U190 (.IN1(enc_round_nr[2]), .IN2(encdec), .IN3(dec_round_nr[2]), .IN4(n43), .Q(
          muxed_round_nr[2]));
   AO22X1 U191 (.IN1(enc_round_nr[1]), .IN2(encdec), .IN3(dec_round_nr[1]), .IN4(n43), .Q(
          muxed_round_nr[1]));
   AO22X1 U192 (.IN1(enc_round_nr[0]), .IN2(encdec), .IN3(dec_round_nr[0]), .IN4(n43), .Q(
          muxed_round_nr[0]));
   aes_encipher_block_test_1 enc_block (.clk(clk), .reset_n(n45), .next(enc_next), .keylen(
          keylen), .round(enc_round_nr), .round_key(round_key), .sboxw(enc_sboxw), .
          new_sboxw(new_sboxw), .block(block), .new_block(enc_new_block), .ready(enc_ready)
          , .test_si(n57), .test_so(n56), .test_se(test_se));
   aes_decipher_block_test_1 dec_block (.clk(clk), .reset_n(n45), .next(dec_next), .keylen(
          keylen), .round(dec_round_nr), .round_key(round_key), .block(block), .new_block(
          dec_new_block), .ready(dec_ready), .test_si(n6), .test_so(n57), .test_se(test_se)
          );
   aes_key_mem_test_1 keymem (.clk(clk), .reset_n(n45), .key(key), .keylen(keylen), .init(
          init), .round(muxed_round_nr), .round_key(round_key), .ready(key_ready), .sboxw(
          keymem_sboxw), .new_sboxw(new_sboxw), .test_si3(test_si3), .test_si2(test_si2), .
          test_si1(n56), .test_so3(n53), .test_so2(test_so2), .test_so1(test_so1), .
          test_se(test_se));
   aes_sbox sbox_inst (.sboxw(muxed_sboxw), .new_sboxw(new_sboxw));
   SDFFARX1 \aes_core_ctrl_reg_reg[1]  (.D(n25), .SI(n9), .SE(test_se), .CLK(clk), .RSTB(
          n45), .Q(aes_core_ctrl_reg[1]), .QN(n6));
   INVX0 U7 (.INP(n46), .ZN(n45));
   NBUFFX2 U8 (.INP(n35), .Z(n11));
   NBUFFX2 U9 (.INP(n33), .Z(n30));
   NBUFFX2 U10 (.INP(n33), .Z(n31));
   NBUFFX2 U11 (.INP(n35), .Z(n22));
   NBUFFX2 U12 (.INP(n33), .Z(n32));
   NBUFFX2 U13 (.INP(n34), .Z(n29));
   NBUFFX2 U14 (.INP(n34), .Z(n27));
   NBUFFX2 U15 (.INP(n34), .Z(n28));
   NBUFFX2 U16 (.INP(n34), .Z(n35));
   NBUFFX2 U17 (.INP(encdec), .Z(n33));
   NBUFFX2 U18 (.INP(encdec), .Z(n34));
   INVX0 U19 (.INP(reset_n), .ZN(n46));
   AO22X1 U150 (.IN1(keymem_sboxw[19]), .IN2(n42), .IN3(enc_sboxw[19]), .IN4(n5), .Q(
          muxed_sboxw[19]));
   AO22X1 U154 (.IN1(keymem_sboxw[17]), .IN2(n42), .IN3(enc_sboxw[17]), .IN4(n7), .Q(
          muxed_sboxw[17]));
   AO22X1 U155 (.IN1(keymem_sboxw[22]), .IN2(n42), .IN3(enc_sboxw[22]), .IN4(n5), .Q(
          muxed_sboxw[22]));
   NOR2X0 U161 (.IN1(n36), .IN2(n49), .QN(enc_next));
   AO22X1 U167 (.IN1(keymem_sboxw[29]), .IN2(n10), .IN3(enc_sboxw[29]), .IN4(n8), .Q(
          muxed_sboxw[29]));
   AO22X1 U174 (.IN1(keymem_sboxw[13]), .IN2(n10), .IN3(enc_sboxw[13]), .IN4(n8), .Q(
          muxed_sboxw[13]));
   AO22X1 U178 (.IN1(keymem_sboxw[5]), .IN2(n10), .IN3(enc_sboxw[5]), .IN4(n8), .Q(
          muxed_sboxw[5]));
   AND3X1 U180 (.IN1(n19), .IN2(n13), .IN3(n20), .Q(n12));
   NAND3X0 U184 (.IN1(n21), .IN2(n9), .IN3(aes_core_ctrl_reg[1]), .QN(n13));
   NOR2X0 U193 (.IN1(init), .IN2(n16), .QN(n17));
   NAND2X1 U194 (.IN1(ready), .IN2(n16), .QN(n15));
   INVX0 U195 (.INP(next), .ZN(n49));
   INVX0 U196 (.INP(n13), .ZN(n47));
   INVX0 U197 (.INP(n42), .ZN(n5));
   INVX0 U198 (.INP(n10), .ZN(n7));
   AO22X1 U199 (.IN1(n16), .IN2(aes_core_ctrl_reg[1]), .IN3(n17), .IN4(n18), .Q(n25));
   OA21X1 U200 (.IN1(n9), .IN2(aes_core_ctrl_reg[1]), .IN3(n19), .Q(n8));
   INVX0 U201 (.INP(n19), .ZN(n48));
   NAND2X0 U202 (.IN1(next), .IN2(n18), .QN(n20));
   INVX0 U203 (.INP(n33), .ZN(n41));
   INVX0 U204 (.INP(n33), .ZN(n38));
   INVX0 U205 (.INP(n33), .ZN(n37));
   INVX0 U206 (.INP(n33), .ZN(n40));
   INVX0 U207 (.INP(n33), .ZN(n39));
   INVX0 U208 (.INP(n34), .ZN(n36));
   INVX0 U209 (.INP(n8), .ZN(n10));
   INVX0 U210 (.INP(n34), .ZN(n44));
   INVX0 U211 (.INP(encdec), .ZN(n43));
   NOR2X0 U212 (.IN1(n11), .IN2(n49), .QN(dec_next));
   INVX0 U213 (.INP(n8), .ZN(n42));
   NOR2X0 U214 (.IN1(aes_core_ctrl_reg[0]), .IN2(aes_core_ctrl_reg[1]), .QN(n18));
   NAND2X0 U215 (.IN1(init), .IN2(n18), .QN(n19));
endmodule

module aes_DW01_add_width3 (A, B, CI, SUM, CO);
input CI;
input [2:0] A;
input [2:0] B;
output CO;
output [2:0] SUM;
wire n4, n5;
   NAND2X2 U1 (.IN1(B[0]), .IN2(A[0]), .QN(n5));
   XNOR2X1 U2 (.IN1(n4), .IN2(A[2]), .Q(SUM[2]));
   NAND3X0 U3 (.IN1(A[1]), .IN2(A[0]), .IN3(B[0]), .QN(n4));
   XNOR2X1 U4 (.IN1(A[1]), .IN2(n5), .Q(SUM[1]));
   XOR2X1 U5 (.IN1(B[0]), .IN2(A[0]), .Q(SUM[0]));
endmodule

module aes_DFT_cntr_scnto_width3_count_to5_rst_mode0_dcod_mode0_0_0 (clk, rst_n, enable, 
       load_n, tercnt_n, count);
input clk, rst_n, enable, load_n;
output tercnt_n;
output [2:0] count;
wire n6, n10, n9, n8, n13, n11, n14, n1;
   aes_DW01_add_width3 add_124 (.A(count), .B({1'b0, 1'b0, enable}), .CI(1'b0), .SUM({n10
          , n9, n8}));
   DFFARX1 \count_int_reg[0]  (.D(n11), .CLK(clk), .RSTB(rst_n), .Q(count[0]));
   DFFARX1 \count_int_reg[1]  (.D(n14), .CLK(clk), .RSTB(rst_n), .Q(count[1]));
   DFFARX1 \count_int_reg[2]  (.D(n13), .CLK(clk), .RSTB(rst_n), .Q(count[2]));
   DFFARX1 tercnt_n_reg_reg (.D(n6), .CLK(clk), .RSTB(rst_n), .QN(tercnt_n));
   INVX1 U4 (.INP(n9), .ZN(n1));
   AND3X1 U5 (.IN1(n8), .IN2(n1), .IN3(n13), .Q(n6));
   AND2X1 U6 (.IN1(load_n), .IN2(n9), .Q(n14));
   AND2X1 U7 (.IN1(n10), .IN2(load_n), .Q(n13));
   AND2X1 U8 (.IN1(load_n), .IN2(n8), .Q(n11));
endmodule

module aes_DFT_decode_width4_0_0 (A, B);
input [2:0] A;
output [7:0] B;
wire n1, n2, n3;
   INVX1 U2 (.INP(A[2]), .ZN(n1));
   INVX1 U3 (.INP(A[1]), .ZN(n2));
   INVX1 U4 (.INP(A[0]), .ZN(n3));
   AND3X1 U5 (.IN1(A[1]), .IN2(A[0]), .IN3(A[2]), .Q(B[7]));
   NOR3X0 U6 (.IN1(n1), .IN2(A[0]), .IN3(n2), .QN(B[6]));
   NOR3X0 U7 (.IN1(n1), .IN2(A[1]), .IN3(n3), .QN(B[5]));
   NOR3X0 U8 (.IN1(n1), .IN2(A[1]), .IN3(A[0]), .QN(B[4]));
   NOR3X0 U9 (.IN1(n2), .IN2(A[2]), .IN3(n3), .QN(B[3]));
   NOR3X0 U10 (.IN1(n2), .IN2(A[2]), .IN3(A[0]), .QN(B[2]));
   NOR3X0 U11 (.IN1(n3), .IN2(A[2]), .IN3(A[1]), .QN(B[1]));
   NOR3X0 U12 (.IN1(A[0]), .IN2(A[2]), .IN3(A[1]), .QN(B[0]));
endmodule

module aes_DFT_or_gate_width4_0_0 (a, b);
input [3:0] a;
output b;
   OR4X1 U1 (.IN1(a[1]), .IN2(a[0]), .IN3(a[3]), .IN4(a[2]), .Q(b));
endmodule

module aes_DFT_clk_control_0_0 (reset, scan_en, clk_enable, fast_clk, slow_clk, 
       fast_clk_enable, slow_clk_enable);
input reset, scan_en, fast_clk, slow_clk;
input [3:0] clk_enable;
output fast_clk_enable, slow_clk_enable;
wire n5, n6, n10, n9, n8, n7, n15, n14, n13, n12, n21, n20, n19, n22, n23, n25, n26, n28, 
       n29, n31, n1, n2, n3, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
       SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
   aes_DFT_cntr_scnto_width3_count_to5_rst_mode0_dcod_mode0_0_0 U_cycle_ctr_i
          (.clk(fast_clk), .rst_n(n2), .enable(n22), .load_n(n25), .tercnt_n(n23), .count({
          n21, n20, n19}));
   aes_DFT_decode_width4_0_0 U_decode_i (.A({n21, n20, n19}), .B({SYNOPSYS_UNCONNECTED__0
          , SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, n15, n14, n13, n12, 
          SYNOPSYS_UNCONNECTED__3}));
   aes_DFT_or_gate_width4_0_0 U_or_tree_i (.a({n10, n9, n8, n7}), .b(n6));
   DFFARX1 pipeline_or_tree_l_reg (.D(n6), .CLK(fast_clk), .RSTB(n2), .Q(n5));
   DFFNARX1 fast_clk_enable_l_reg (.D(n31), .CLK(fast_clk), .RSTB(n2), .Q(fast_clk_enable)
          );
   DFFNARX1 slow_clk_enable_l_reg (.D(n29), .CLK(slow_clk), .RSTB(n2), .Q(slow_clk_enable)
          , .QN(n1));
   DFFARX1 load_n_meta_0_l_reg (.D(n1), .CLK(fast_clk), .RSTB(n2), .Q(n28));
   DFFARX1 load_n_meta_1_l_reg (.D(n28), .CLK(fast_clk), .RSTB(n2), .Q(n26));
   DFFARX1 load_n_meta_2_l_reg (.D(n26), .CLK(fast_clk), .RSTB(n2), .Q(n25));
   NOR2X2 U3 (.IN1(fast_clk_enable), .IN2(n3), .QN(n29));
   INVX1 U4 (.INP(reset), .ZN(n2));
   INVX1 U5 (.INP(scan_en), .ZN(n3));
   AND2X1 U6 (.IN1(n14), .IN2(clk_enable[2]), .Q(n9));
   AND2X1 U7 (.IN1(n13), .IN2(clk_enable[1]), .Q(n8));
   AND2X1 U8 (.IN1(n12), .IN2(clk_enable[0]), .Q(n7));
   AND3X1 U9 (.IN1(n3), .IN2(n1), .IN3(n5), .Q(n31));
   AND2X1 U10 (.IN1(n23), .IN2(n3), .Q(n22));
   AND2X1 U11 (.IN1(n15), .IN2(clk_enable[3]), .Q(n10));
endmodule

module aes_DFT_gf_mux_0_0 (fast_clk_enable, slow_clk_enable, pll_bypass, test_mode, 
       scan_en, fast_gate, slow_gate);
input fast_clk_enable, slow_clk_enable, pll_bypass, test_mode, scan_en;
output fast_gate, slow_gate;
wire n1, n2;
   OA21X2 U1 (.IN1(n2), .IN2(pll_bypass), .IN3(test_mode), .Q(slow_gate));
   INVX1 U2 (.INP(fast_clk_enable), .ZN(n1));
   AND2X1 U3 (.IN1(slow_clk_enable), .IN2(scan_en), .Q(n2));
   OAI21X1 U4 (.IN1(n1), .IN2(pll_bypass), .IN3(test_mode), .QN(fast_gate));
endmodule

module aes_mselector_n2_m1_0 (DATA1_0, DATA2_0, CONTROL1, CONTROL2, Z_0);
input DATA1_0, DATA2_0, CONTROL1, CONTROL2;
output Z_0;
   AO22X1 U2 (.IN1(DATA2_0), .IN2(CONTROL2), .IN3(DATA1_0), .IN4(CONTROL1), .Q(Z_0));
endmodule

module aes_mselector_n2_m1 (DATA1_0, DATA2_0, CONTROL1, CONTROL2, Z_0);
input DATA1_0, DATA2_0, CONTROL1, CONTROL2;
output Z_0;
   AO22X1 U2 (.IN1(DATA2_0), .IN2(CONTROL2), .IN3(DATA1_0), .IN4(CONTROL1), .Q(Z_0));
endmodule

module aes_DFT_clk_mux_0 (fast_clk, scan_en, test_mode, reset, pll_bypass, slow_clk, 
       clk_enable, clk);
input fast_clk, scan_en, test_mode, reset, pll_bypass, slow_clk;
input [3:0] clk_enable;
output clk;
wire n6, n7, n21, n23, n2, n3, n4;
   aes_DFT_clk_control_0_0 U_clk_control_i_0 (.reset(reset), .scan_en(scan_en), .
          clk_enable(clk_enable), .fast_clk(fast_clk), .slow_clk(slow_clk), .
          fast_clk_enable(n7), .slow_clk_enable(n6));
   aes_DFT_gf_mux_0_0 U_gf_mux_0 (.fast_clk_enable(n7), .slow_clk_enable(n6), .pll_bypass(
          pll_bypass), .test_mode(test_mode), .scan_en(scan_en), .fast_gate(n23), .
          slow_gate(n21));
   aes_mselector_n2_m1_0 U2 (.DATA1_0(fast_clk), .DATA2_0(n2), .CONTROL1(n23), .CONTROL2(
          n4), .Z_0(clk));
   aes_mselector_n2_m1 U3 (.DATA1_0(slow_clk), .DATA2_0(1'b0), .CONTROL1(n21), .CONTROL2(
          n3), .Z_0(n2));
   INVX1 U5 (.INP(n21), .ZN(n3));
   INVX1 U6 (.INP(n23), .ZN(n4));
endmodule

module aes_DFT_clk_chain_0 (clk, se, si, so, clk_ctrl_data);
input clk, se, si;
output so;
output [3:0] clk_ctrl_data;
wire n7, n14, n21, n28, n1;
   assign clk_ctrl_data[3] = so;
   DFFNX1 \U_shftreg_0/ff_3/q_reg  (.D(n28), .CLK(clk), .Q(clk_ctrl_data[0]));
   DFFNX1 \U_shftreg_0/ff_2/q_reg  (.D(n21), .CLK(clk), .Q(clk_ctrl_data[1]));
   DFFNX1 \U_shftreg_0/ff_1/q_reg  (.D(n14), .CLK(clk), .Q(clk_ctrl_data[2]));
   DFFNX1 \U_shftreg_0/ff_0/q_reg  (.D(n7), .CLK(clk), .Q(so));
   INVX1 U1 (.INP(se), .ZN(n1));
   AO22X1 U2 (.IN1(so), .IN2(n1), .IN3(se), .IN4(clk_ctrl_data[2]), .Q(n7));
   AO22X1 U3 (.IN1(si), .IN2(se), .IN3(clk_ctrl_data[0]), .IN4(n1), .Q(n28));
   AO22X1 U4 (.IN1(clk_ctrl_data[0]), .IN2(se), .IN3(clk_ctrl_data[1]), .IN4(n1), .Q(n21)
          );
   AO22X1 U5 (.IN1(clk_ctrl_data[2]), .IN2(n1), .IN3(clk_ctrl_data[1]), .IN4(se), .Q(n14)
          );
endmodule

module aes (clk, TEST_SE, TEST_SI1, TEST_SI2, TEST_SI3, reset_n, cs, we, address, 
       write_data, read_data, TEST_SO1, TEST_SO2, TEST_SO3, scan_clk, SCAN_MODE, 
       internal_pll_bypass, pll_bypass, pll_reset, test_si4, test_so4);
input clk, TEST_SE, TEST_SI1, TEST_SI2, TEST_SI3, reset_n, cs, we, scan_clk, SCAN_MODE, 
       internal_pll_bypass, pll_bypass, pll_reset, test_si4;
input [7:0] address;
input [31:0] write_data;
output TEST_SO1, TEST_SO2, TEST_SO3, test_so4;
output [31:0] read_data;
wire n1562, core_init, core_next, core_encdec, core_keylen, core_ready, core_valid, 
       valid_reg, ready_reg, init_new, next_new, N62, N64, N108, N109, n552, n555, n556, 
       n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570
       , n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
       n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597
       , n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
       n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624
       , n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, 
       n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651
       , n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
       n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678
       , n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
       n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705
       , n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
       n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732
       , n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
       n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759
       , n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, 
       n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786
       , n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
       n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813
       , n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, 
       n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840
       , n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, 
       n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867
       , n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, 
       n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894
       , n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
       n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921
       , n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, 
       n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948
       , n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
       n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975
       , n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, 
       n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, 
       n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013
       , n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, 
       n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036
       , n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, 
       n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059
       , n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, 
       n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082
       , n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
       n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105
       , n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, 
       n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128
       , n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
       n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151
       , n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
       \clk_ctrl_data[0] , \clk_ctrl_data[1] , \clk_ctrl_data[2] , \clk_ctrl_data[3] , 
       n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173
       , n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
       n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196
       , n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, 
       n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219
       , n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, 
       n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242
       , n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, 
       n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265
       , n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, 
       n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288
       , n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
       n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311
       , n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
       n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334
       , n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
       n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357
       , n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
       n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380
       , n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, 
       n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403
       , n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
       n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1429, n1430, n1431, n1432
       , n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
       n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455
       , n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, 
       n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478
       , n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
       n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501
       , n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
       n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524
       , n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
       n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547
       , n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1560, 
       TEST_SE_buf_net0, TEST_SE_buf_net1, n1562_buf_net0, n1562_buf_net1;
wire [255:0] core_key;
wire [127:0] core_block;
wire [127:0] core_result;
wire [127:0] result_reg;
   assign test_so4 = valid_reg;
   SDFFARX1 \key_reg_reg[0][31]  (.D(n1013), .SI(n1389), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[255]), .QN(n1388));
   SDFFARX1 \key_reg_reg[0][30]  (.D(n1012), .SI(n1390), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[254]), .QN(n1389));
   SDFFARX1 \key_reg_reg[0][29]  (.D(n1011), .SI(n1391), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[253]), .QN(n1390));
   SDFFARX1 \key_reg_reg[0][28]  (.D(n1010), .SI(n1392), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[252]), .QN(n1391));
   SDFFARX1 \key_reg_reg[0][27]  (.D(n1009), .SI(n1393), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[251]), .QN(n1392));
   SDFFARX1 \key_reg_reg[0][26]  (.D(n1008), .SI(n1394), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[250]), .QN(n1393));
   SDFFARX1 \key_reg_reg[0][25]  (.D(n1007), .SI(n1395), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[249]), .QN(n1394));
   SDFFARX1 \key_reg_reg[0][24]  (.D(n1006), .SI(n1396), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[248]), .QN(n1395));
   SDFFARX1 \key_reg_reg[0][23]  (.D(n1005), .SI(n1397), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[247]), .QN(n1396));
   SDFFARX1 \key_reg_reg[0][22]  (.D(n1004), .SI(n1398), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[246]), .QN(n1397));
   SDFFARX1 \key_reg_reg[0][21]  (.D(n1003), .SI(n1399), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[245]), .QN(n1398));
   SDFFARX1 \key_reg_reg[0][20]  (.D(n1002), .SI(n1400), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[244]), .QN(n1399));
   SDFFARX1 \key_reg_reg[0][19]  (.D(n1001), .SI(n1401), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[243]), .QN(n1400));
   SDFFARX1 \key_reg_reg[0][18]  (.D(n1000), .SI(n1402), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[242]), .QN(n1401));
   SDFFARX1 \key_reg_reg[0][17]  (.D(n999), .SI(n1403), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[241]), .QN(n1402));
   SDFFARX1 \key_reg_reg[0][16]  (.D(n998), .SI(n1404), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[240]), .QN(n1403));
   SDFFARX1 \key_reg_reg[0][15]  (.D(n997), .SI(n1405), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[239]), .QN(n1404));
   SDFFARX1 \key_reg_reg[0][14]  (.D(n996), .SI(n1406), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[238]), .QN(n1405));
   SDFFARX1 \key_reg_reg[0][13]  (.D(n995), .SI(n1407), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[237]), .QN(n1406));
   SDFFARX1 \key_reg_reg[0][12]  (.D(n994), .SI(n1408), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[236]), .QN(n1407));
   SDFFARX1 \key_reg_reg[0][11]  (.D(n993), .SI(n1409), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[235]), .QN(n1408));
   SDFFARX1 \key_reg_reg[0][10]  (.D(n992), .SI(n1410), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[234]), .QN(n1409));
   SDFFARX1 \key_reg_reg[0][9]  (.D(n991), .SI(n1411), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[233]), .QN(n1410));
   SDFFARX1 \key_reg_reg[0][8]  (.D(n990), .SI(n1412), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[232]), .QN(n1411));
   SDFFARX1 \key_reg_reg[0][7]  (.D(n989), .SI(n1413), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[231]), .QN(n1412));
   SDFFARX1 \key_reg_reg[0][6]  (.D(n988), .SI(n1414), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[230]), .QN(n1413));
   SDFFARX1 \key_reg_reg[0][5]  (.D(n987), .SI(n1415), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[229]), .QN(n1414));
   SDFFARX1 \key_reg_reg[0][4]  (.D(n986), .SI(n1416), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[228]), .QN(n1415));
   SDFFARX1 \key_reg_reg[0][3]  (.D(n985), .SI(n1417), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[227]), .QN(n1416));
   SDFFARX1 \key_reg_reg[0][2]  (.D(n984), .SI(n1418), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[226]), .QN(n1417));
   SDFFARX1 \key_reg_reg[0][1]  (.D(n983), .SI(n1419), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[225]), .QN(n1418));
   SDFFARX1 \key_reg_reg[0][0]  (.D(n982), .SI(n1420), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[224]), .QN(n1419));
   SDFFARX1 \key_reg_reg[1][31]  (.D(n981), .SI(n1357), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[223]), .QN(n1356));
   SDFFARX1 \key_reg_reg[1][30]  (.D(n980), .SI(n1358), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1143), .Q(core_key[222]), .QN(n1357));
   SDFFARX1 \key_reg_reg[1][29]  (.D(n979), .SI(n1359), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1144), .Q(core_key[221]), .QN(n1358));
   SDFFARX1 \key_reg_reg[1][28]  (.D(n978), .SI(n1360), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1145), .Q(core_key[220]), .QN(n1359));
   SDFFARX1 \key_reg_reg[1][27]  (.D(n977), .SI(n1361), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1092), .Q(core_key[219]), .QN(n1360));
   SDFFARX1 \key_reg_reg[1][26]  (.D(n976), .SI(n1362), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1103), .Q(core_key[218]), .QN(n1361));
   SDFFARX1 \key_reg_reg[1][25]  (.D(n975), .SI(n1363), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1106), .Q(core_key[217]), .QN(n1362));
   SDFFARX1 \key_reg_reg[1][24]  (.D(n974), .SI(n1364), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1089), .Q(core_key[216]), .QN(n1363));
   SDFFARX1 \key_reg_reg[1][23]  (.D(n973), .SI(n1365), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1077), .Q(core_key[215]), .QN(n1364));
   SDFFARX1 \key_reg_reg[1][22]  (.D(n972), .SI(n1366), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1076), .Q(core_key[214]), .QN(n1365));
   SDFFARX1 \key_reg_reg[1][21]  (.D(n971), .SI(n1367), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1075), .Q(core_key[213]), .QN(n1366));
   SDFFARX1 \key_reg_reg[1][20]  (.D(n970), .SI(n1368), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1078), .Q(core_key[212]), .QN(n1367));
   SDFFARX1 \key_reg_reg[1][19]  (.D(n969), .SI(n1369), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1091), .Q(core_key[211]), .QN(n1368));
   SDFFARX1 \key_reg_reg[1][18]  (.D(n968), .SI(n1370), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1090), .Q(core_key[210]), .QN(n1369));
   SDFFARX1 \key_reg_reg[1][17]  (.D(n967), .SI(n1371), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1105), .Q(core_key[209]), .QN(n1370));
   SDFFARX1 \key_reg_reg[1][16]  (.D(n966), .SI(n1372), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1104), .Q(core_key[208]), .QN(n1371));
   SDFFARX1 \key_reg_reg[1][15]  (.D(n965), .SI(n1373), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1092), .Q(core_key[207]), .QN(n1372));
   SDFFARX1 \key_reg_reg[1][14]  (.D(n964), .SI(n1374), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1103), .Q(core_key[206]), .QN(n1373));
   SDFFARX1 \key_reg_reg[1][13]  (.D(n963), .SI(n1375), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1106), .Q(core_key[205]), .QN(n1374));
   SDFFARX1 \key_reg_reg[1][12]  (.D(n962), .SI(n1376), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1089), .Q(core_key[204]), .QN(n1375));
   SDFFARX1 \key_reg_reg[1][11]  (.D(n961), .SI(n1377), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[203]), .QN(n1376));
   SDFFARX1 \key_reg_reg[1][10]  (.D(n960), .SI(n1378), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[202]), .QN(n1377));
   SDFFARX1 \key_reg_reg[1][9]  (.D(n959), .SI(n1379), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[201]), .QN(n1378));
   SDFFARX1 \key_reg_reg[1][8]  (.D(n958), .SI(n1380), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[200]), .QN(n1379));
   SDFFARX1 \key_reg_reg[1][7]  (.D(n957), .SI(n1381), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[199]), .QN(n1380));
   SDFFARX1 \key_reg_reg[1][6]  (.D(n956), .SI(n1382), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[198]), .QN(n1381));
   SDFFARX1 \key_reg_reg[1][5]  (.D(n955), .SI(n1383), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[197]), .QN(n1382));
   SDFFARX1 \key_reg_reg[1][4]  (.D(n954), .SI(n1384), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[196]), .QN(n1383));
   SDFFARX1 \key_reg_reg[1][3]  (.D(n953), .SI(n1385), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[195]), .QN(n1384));
   SDFFARX1 \key_reg_reg[1][2]  (.D(n952), .SI(n1386), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[194]), .QN(n1385));
   SDFFARX1 \key_reg_reg[1][1]  (.D(n951), .SI(n1387), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[193]), .QN(n1386));
   SDFFARX1 \key_reg_reg[1][0]  (.D(n950), .SI(n1388), .SE(TEST_SE), .CLK(n1562), .RSTB(
          reset_n), .Q(core_key[192]), .QN(n1387));
   SDFFARX1 \key_reg_reg[2][31]  (.D(n949), .SI(n1325), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[191]), .QN(n1324));
   SDFFARX1 \key_reg_reg[2][30]  (.D(n948), .SI(n1326), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[190]), .QN(n1325));
   SDFFARX1 \key_reg_reg[2][29]  (.D(n947), .SI(n1327), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[189]), .QN(n1326));
   SDFFARX1 \key_reg_reg[2][28]  (.D(n946), .SI(n1328), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[188]), .QN(n1327));
   SDFFARX1 \key_reg_reg[2][27]  (.D(n945), .SI(n1329), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[187]), .QN(n1328));
   SDFFARX1 \key_reg_reg[2][26]  (.D(n944), .SI(n1330), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[186]), .QN(n1329));
   SDFFARX1 \key_reg_reg[2][25]  (.D(n943), .SI(n1331), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[185]), .QN(n1330));
   SDFFARX1 \key_reg_reg[2][24]  (.D(n942), .SI(n1332), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[184]), .QN(n1331));
   SDFFARX1 \key_reg_reg[2][23]  (.D(n941), .SI(n1333), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[183]), .QN(n1332));
   SDFFARX1 \key_reg_reg[2][22]  (.D(n940), .SI(n1334), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[182]), .QN(n1333));
   SDFFARX1 \key_reg_reg[2][21]  (.D(n939), .SI(n1335), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[181]), .QN(n1334));
   SDFFARX1 \key_reg_reg[2][20]  (.D(n938), .SI(n1336), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[180]), .QN(n1335));
   SDFFARX1 \key_reg_reg[2][19]  (.D(n937), .SI(n1337), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1102), .Q(core_key[179]), .QN(n1336));
   SDFFARX1 \key_reg_reg[2][18]  (.D(n936), .SI(n1338), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[178]), .QN(n1337));
   SDFFARX1 \key_reg_reg[2][17]  (.D(n935), .SI(n1339), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[177]), .QN(n1338));
   SDFFARX1 \key_reg_reg[2][16]  (.D(n934), .SI(n1340), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[176]), .QN(n1339));
   SDFFARX1 \key_reg_reg[2][15]  (.D(n933), .SI(n1341), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[175]), .QN(n1340));
   SDFFARX1 \key_reg_reg[2][14]  (.D(n932), .SI(n1342), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[174]), .QN(n1341));
   SDFFARX1 \key_reg_reg[2][13]  (.D(n931), .SI(n1343), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[173]), .QN(n1342));
   SDFFARX1 \key_reg_reg[2][12]  (.D(n930), .SI(n1344), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[172]), .QN(n1343));
   SDFFARX1 \key_reg_reg[2][11]  (.D(n929), .SI(n1345), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[171]), .QN(n1344));
   SDFFARX1 \key_reg_reg[2][10]  (.D(n928), .SI(n1346), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[170]), .QN(n1345));
   SDFFARX1 \key_reg_reg[2][9]  (.D(n927), .SI(n1347), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[169]), .QN(n1346));
   SDFFARX1 \key_reg_reg[2][8]  (.D(n926), .SI(n1348), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[168]), .QN(n1347));
   SDFFARX1 \key_reg_reg[2][7]  (.D(n925), .SI(n1349), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1101), .Q(core_key[167]), .QN(n1348));
   SDFFARX1 \key_reg_reg[2][6]  (.D(n924), .SI(n1350), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[166]), .QN(n1349));
   SDFFARX1 \key_reg_reg[2][5]  (.D(n923), .SI(n1351), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[165]), .QN(n1350));
   SDFFARX1 \key_reg_reg[2][4]  (.D(n922), .SI(n1352), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[164]), .QN(n1351));
   SDFFARX1 \key_reg_reg[2][3]  (.D(n921), .SI(n1353), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[163]), .QN(n1352));
   SDFFARX1 \key_reg_reg[2][2]  (.D(n920), .SI(n1354), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[162]), .QN(n1353));
   SDFFARX1 \key_reg_reg[2][1]  (.D(n919), .SI(n1355), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[161]), .QN(n1354));
   SDFFARX1 \key_reg_reg[2][0]  (.D(n918), .SI(n1356), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[160]), .QN(n1355));
   SDFFARX1 \key_reg_reg[3][31]  (.D(n917), .SI(n1293), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[159]), .QN(n1292));
   SDFFARX1 \key_reg_reg[3][30]  (.D(n916), .SI(n1294), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[158]), .QN(n1293));
   SDFFARX1 \key_reg_reg[3][29]  (.D(n915), .SI(n1295), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[157]), .QN(n1294));
   SDFFARX1 \key_reg_reg[3][28]  (.D(n914), .SI(n1296), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[156]), .QN(n1295));
   SDFFARX1 \key_reg_reg[3][27]  (.D(n913), .SI(n1297), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1100), .Q(core_key[155]), .QN(n1296));
   SDFFARX1 \key_reg_reg[3][26]  (.D(n912), .SI(n1298), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[154]), .QN(n1297));
   SDFFARX1 \key_reg_reg[3][25]  (.D(n911), .SI(n1299), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[153]), .QN(n1298));
   SDFFARX1 \key_reg_reg[3][24]  (.D(n910), .SI(n1300), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[152]), .QN(n1299));
   SDFFARX1 \key_reg_reg[3][23]  (.D(n909), .SI(n1301), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[151]), .QN(n1300));
   SDFFARX1 \key_reg_reg[3][22]  (.D(n908), .SI(n1302), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[150]), .QN(n1301));
   SDFFARX1 \key_reg_reg[3][21]  (.D(n907), .SI(n1303), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[149]), .QN(n1302));
   SDFFARX1 \key_reg_reg[3][20]  (.D(n906), .SI(n1304), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[148]), .QN(n1303));
   SDFFARX1 \key_reg_reg[3][19]  (.D(n905), .SI(n1305), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[147]), .QN(n1304));
   SDFFARX1 \key_reg_reg[3][18]  (.D(n904), .SI(n1306), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[146]), .QN(n1305));
   SDFFARX1 \key_reg_reg[3][17]  (.D(n903), .SI(n1307), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[145]), .QN(n1306));
   SDFFARX1 \key_reg_reg[3][16]  (.D(n902), .SI(n1308), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[144]), .QN(n1307));
   SDFFARX1 \key_reg_reg[3][15]  (.D(n901), .SI(n1309), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1099), .Q(core_key[143]), .QN(n1308));
   SDFFARX1 \key_reg_reg[3][14]  (.D(n900), .SI(n1310), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[142]), .QN(n1309));
   SDFFARX1 \key_reg_reg[3][13]  (.D(n899), .SI(n1311), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[141]), .QN(n1310));
   SDFFARX1 \key_reg_reg[3][12]  (.D(n898), .SI(n1312), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[140]), .QN(n1311));
   SDFFARX1 \key_reg_reg[3][11]  (.D(n897), .SI(n1313), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[139]), .QN(n1312));
   SDFFARX1 \key_reg_reg[3][10]  (.D(n896), .SI(n1314), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[138]), .QN(n1313));
   SDFFARX1 \key_reg_reg[3][9]  (.D(n895), .SI(n1315), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[137]), .QN(n1314));
   SDFFARX1 \key_reg_reg[3][8]  (.D(n894), .SI(n1316), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[136]), .QN(n1315));
   SDFFARX1 \key_reg_reg[3][7]  (.D(n893), .SI(n1317), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[135]), .QN(n1316));
   SDFFARX1 \key_reg_reg[3][6]  (.D(n892), .SI(n1318), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[134]), .QN(n1317));
   SDFFARX1 \key_reg_reg[3][5]  (.D(n891), .SI(n1319), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[133]), .QN(n1318));
   SDFFARX1 \key_reg_reg[3][4]  (.D(n890), .SI(n1320), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[132]), .QN(n1319));
   SDFFARX1 \key_reg_reg[3][3]  (.D(n889), .SI(n1321), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1098), .Q(core_key[131]), .QN(n1320));
   SDFFARX1 \key_reg_reg[3][2]  (.D(n888), .SI(n1322), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[130]), .QN(n1321));
   SDFFARX1 \key_reg_reg[3][1]  (.D(n887), .SI(n1323), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[129]), .QN(n1322));
   SDFFARX1 \key_reg_reg[3][0]  (.D(n886), .SI(n1324), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[128]), .QN(n1323));
   SDFFARX1 \key_reg_reg[4][31]  (.D(n885), .SI(n1261), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[127]), .QN(n1260));
   SDFFARX1 \key_reg_reg[4][30]  (.D(n884), .SI(n1262), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[126]), .QN(n1261));
   SDFFARX1 \key_reg_reg[4][29]  (.D(n883), .SI(n1263), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[125]), .QN(n1262));
   SDFFARX1 \key_reg_reg[4][28]  (.D(n882), .SI(n1264), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[124]), .QN(n1263));
   SDFFARX1 \key_reg_reg[4][27]  (.D(n881), .SI(n1265), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[123]), .QN(n1264));
   SDFFARX1 \key_reg_reg[4][26]  (.D(n880), .SI(n1266), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[122]), .QN(n1265));
   SDFFARX1 \key_reg_reg[4][25]  (.D(n879), .SI(n1267), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[121]), .QN(n1266));
   SDFFARX1 \key_reg_reg[4][24]  (.D(n878), .SI(n1268), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[120]), .QN(n1267));
   SDFFARX1 \key_reg_reg[4][23]  (.D(n877), .SI(n1269), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1097), .Q(core_key[119]), .QN(n1268));
   SDFFARX1 \key_reg_reg[4][22]  (.D(n876), .SI(n1270), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[118]), .QN(n1269));
   SDFFARX1 \key_reg_reg[4][21]  (.D(n875), .SI(n1271), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[117]), .QN(n1270));
   SDFFARX1 \key_reg_reg[4][20]  (.D(n874), .SI(n1272), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[116]), .QN(n1271));
   SDFFARX1 \key_reg_reg[4][19]  (.D(n873), .SI(n1273), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[115]), .QN(n1272));
   SDFFARX1 \key_reg_reg[4][18]  (.D(n872), .SI(n1274), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[114]), .QN(n1273));
   SDFFARX1 \key_reg_reg[4][17]  (.D(n871), .SI(n1275), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[113]), .QN(n1274));
   SDFFARX1 \key_reg_reg[4][16]  (.D(n870), .SI(n1276), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[112]), .QN(n1275));
   SDFFARX1 \key_reg_reg[4][15]  (.D(n869), .SI(n1277), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[111]), .QN(n1276));
   SDFFARX1 \key_reg_reg[4][14]  (.D(n868), .SI(n1278), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[110]), .QN(n1277));
   SDFFARX1 \key_reg_reg[4][13]  (.D(n867), .SI(n1279), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[109]), .QN(n1278));
   SDFFARX1 \key_reg_reg[4][12]  (.D(n866), .SI(n1280), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[108]), .QN(n1279));
   SDFFARX1 \key_reg_reg[4][11]  (.D(n865), .SI(n1281), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1096), .Q(core_key[107]), .QN(n1280));
   SDFFARX1 \key_reg_reg[4][10]  (.D(n864), .SI(n1282), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[106]), .QN(n1281));
   SDFFARX1 \key_reg_reg[4][9]  (.D(n863), .SI(n1283), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[105]), .QN(n1282));
   SDFFARX1 \key_reg_reg[4][8]  (.D(n862), .SI(n1284), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[104]), .QN(n1283));
   SDFFARX1 \key_reg_reg[4][7]  (.D(n861), .SI(n1285), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[103]), .QN(n1284));
   SDFFARX1 \key_reg_reg[4][6]  (.D(n860), .SI(n1286), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[102]), .QN(n1285));
   SDFFARX1 \key_reg_reg[4][5]  (.D(n859), .SI(n1287), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[101]), .QN(n1286));
   SDFFARX1 \key_reg_reg[4][4]  (.D(n858), .SI(n1288), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[100]), .QN(n1287));
   SDFFARX1 \key_reg_reg[4][3]  (.D(n857), .SI(n1289), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[99]), .QN(n1288));
   SDFFARX1 \key_reg_reg[4][2]  (.D(n856), .SI(n1290), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[98]), .QN(n1289));
   SDFFARX1 \key_reg_reg[4][1]  (.D(n855), .SI(n1291), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[97]), .QN(n1290));
   SDFFARX1 \key_reg_reg[4][0]  (.D(n854), .SI(n1292), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[96]), .QN(n1291));
   SDFFARX1 \key_reg_reg[5][31]  (.D(n853), .SI(n1229), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1095), .Q(core_key[95]), .QN(n1228));
   SDFFARX1 \key_reg_reg[5][30]  (.D(n852), .SI(n1230), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[94]), .QN(n1229));
   SDFFARX1 \key_reg_reg[5][29]  (.D(n851), .SI(n1231), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[93]), .QN(n1230));
   SDFFARX1 \key_reg_reg[5][28]  (.D(n850), .SI(n1232), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[92]), .QN(n1231));
   SDFFARX1 \key_reg_reg[5][27]  (.D(n849), .SI(n1233), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[91]), .QN(n1232));
   SDFFARX1 \key_reg_reg[5][26]  (.D(n848), .SI(n1234), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[90]), .QN(n1233));
   SDFFARX1 \key_reg_reg[5][25]  (.D(n847), .SI(n1235), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[89]), .QN(n1234));
   SDFFARX1 \key_reg_reg[5][24]  (.D(n846), .SI(n1236), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[88]), .QN(n1235));
   SDFFARX1 \key_reg_reg[5][23]  (.D(n845), .SI(n1237), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[87]), .QN(n1236));
   SDFFARX1 \key_reg_reg[5][22]  (.D(n844), .SI(n1238), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[86]), .QN(n1237));
   SDFFARX1 \key_reg_reg[5][21]  (.D(n843), .SI(n1239), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[85]), .QN(n1238));
   SDFFARX1 \key_reg_reg[5][20]  (.D(n842), .SI(n1240), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[84]), .QN(n1239));
   SDFFARX1 \key_reg_reg[5][19]  (.D(n841), .SI(n1241), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1094), .Q(core_key[83]), .QN(n1240));
   SDFFARX1 \key_reg_reg[5][18]  (.D(n840), .SI(n1242), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[82]), .QN(n1241));
   SDFFARX1 \key_reg_reg[5][17]  (.D(n839), .SI(n1243), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[81]), .QN(n1242));
   SDFFARX1 \key_reg_reg[5][16]  (.D(n838), .SI(n1244), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[80]), .QN(n1243));
   SDFFARX1 \key_reg_reg[5][15]  (.D(n837), .SI(n1245), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[79]), .QN(n1244));
   SDFFARX1 \key_reg_reg[5][14]  (.D(n836), .SI(n1246), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[78]), .QN(n1245));
   SDFFARX1 \key_reg_reg[5][13]  (.D(n835), .SI(n1247), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[77]), .QN(n1246));
   SDFFARX1 \key_reg_reg[5][12]  (.D(n834), .SI(n1248), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[76]), .QN(n1247));
   SDFFARX1 \key_reg_reg[5][11]  (.D(n833), .SI(n1249), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[75]), .QN(n1248));
   SDFFARX1 \key_reg_reg[5][10]  (.D(n832), .SI(n1250), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[74]), .QN(n1249));
   SDFFARX1 \key_reg_reg[5][9]  (.D(n831), .SI(n1251), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[73]), .QN(n1250));
   SDFFARX1 \key_reg_reg[5][8]  (.D(n830), .SI(n1252), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[72]), .QN(n1251));
   SDFFARX1 \key_reg_reg[5][7]  (.D(n829), .SI(n1253), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1093), .Q(core_key[71]), .QN(n1252));
   SDFFARX1 \key_reg_reg[5][6]  (.D(n828), .SI(n1254), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1146), .Q(core_key[70]), .QN(n1253));
   SDFFARX1 \key_reg_reg[5][5]  (.D(n827), .SI(n1255), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[69]), .QN(n1254));
   SDFFARX1 \key_reg_reg[5][4]  (.D(n826), .SI(n1256), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[68]), .QN(n1255));
   SDFFARX1 \key_reg_reg[5][3]  (.D(n825), .SI(n1257), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[67]), .QN(n1256));
   SDFFARX1 \key_reg_reg[5][2]  (.D(n824), .SI(n1258), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[66]), .QN(n1257));
   SDFFARX1 \key_reg_reg[5][1]  (.D(n823), .SI(n1259), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[65]), .QN(n1258));
   SDFFARX1 \key_reg_reg[5][0]  (.D(n822), .SI(n1260), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[64]), .QN(n1259));
   SDFFARX1 \key_reg_reg[6][31]  (.D(n821), .SI(n1197), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[63]), .QN(n1196));
   SDFFARX1 \key_reg_reg[6][30]  (.D(n820), .SI(n1198), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[62]), .QN(n1197));
   SDFFARX1 \key_reg_reg[6][29]  (.D(n819), .SI(n1199), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[61]), .QN(n1198));
   SDFFARX1 \key_reg_reg[6][28]  (.D(n818), .SI(n1200), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[60]), .QN(n1199));
   SDFFARX1 \key_reg_reg[6][27]  (.D(n817), .SI(n1201), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[59]), .QN(n1200));
   SDFFARX1 \key_reg_reg[6][26]  (.D(n816), .SI(n1202), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1088), .Q(core_key[58]), .QN(n1201));
   SDFFARX1 \key_reg_reg[6][25]  (.D(n815), .SI(n1203), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[57]), .QN(n1202));
   SDFFARX1 \key_reg_reg[6][24]  (.D(n814), .SI(n1204), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[56]), .QN(n1203));
   SDFFARX1 \key_reg_reg[6][23]  (.D(n813), .SI(n1205), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[55]), .QN(n1204));
   SDFFARX1 \key_reg_reg[6][22]  (.D(n812), .SI(n1206), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[54]), .QN(n1205));
   SDFFARX1 \key_reg_reg[6][21]  (.D(n811), .SI(n1207), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[53]), .QN(n1206));
   SDFFARX1 \key_reg_reg[6][20]  (.D(n810), .SI(n1208), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[52]), .QN(n1207));
   SDFFARX1 \key_reg_reg[6][19]  (.D(n809), .SI(n1209), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[51]), .QN(n1208));
   SDFFARX1 \key_reg_reg[6][18]  (.D(n808), .SI(n1210), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[50]), .QN(n1209));
   SDFFARX1 \key_reg_reg[6][17]  (.D(n807), .SI(n1211), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[49]), .QN(n1210));
   SDFFARX1 \key_reg_reg[6][16]  (.D(n806), .SI(n1212), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[48]), .QN(n1211));
   SDFFARX1 \key_reg_reg[6][15]  (.D(n805), .SI(n1213), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[47]), .QN(n1212));
   SDFFARX1 \key_reg_reg[6][14]  (.D(n804), .SI(n1214), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1087), .Q(core_key[46]), .QN(n1213));
   SDFFARX1 \key_reg_reg[6][13]  (.D(n803), .SI(n1215), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[45]), .QN(n1214));
   SDFFARX1 \key_reg_reg[6][12]  (.D(n802), .SI(n1216), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[44]), .QN(n1215));
   SDFFARX1 \key_reg_reg[6][11]  (.D(n801), .SI(n1217), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[43]), .QN(n1216));
   SDFFARX1 \key_reg_reg[6][10]  (.D(n800), .SI(n1218), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[42]), .QN(n1217));
   SDFFARX1 \key_reg_reg[6][9]  (.D(n799), .SI(n1219), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[41]), .QN(n1218));
   SDFFARX1 \key_reg_reg[6][8]  (.D(n798), .SI(n1220), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[40]), .QN(n1219));
   SDFFARX1 \key_reg_reg[6][7]  (.D(n797), .SI(n1221), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[39]), .QN(n1220));
   SDFFARX1 \key_reg_reg[6][6]  (.D(n796), .SI(n1222), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[38]), .QN(n1221));
   SDFFARX1 \key_reg_reg[6][5]  (.D(n795), .SI(n1223), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[37]), .QN(n1222));
   SDFFARX1 \key_reg_reg[6][4]  (.D(n794), .SI(n1224), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[36]), .QN(n1223));
   SDFFARX1 \key_reg_reg[6][3]  (.D(n793), .SI(n1225), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[35]), .QN(n1224));
   SDFFARX1 \key_reg_reg[6][2]  (.D(n792), .SI(n1226), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1086), .Q(core_key[34]), .QN(n1225));
   SDFFARX1 \key_reg_reg[6][1]  (.D(n791), .SI(n1227), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[33]), .QN(n1226));
   SDFFARX1 \key_reg_reg[6][0]  (.D(n790), .SI(n1228), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[32]), .QN(n1227));
   SDFFARX1 \key_reg_reg[7][31]  (.D(n789), .SI(n1165), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[31]), .QN(n1164));
   SDFFARX1 \key_reg_reg[7][30]  (.D(n788), .SI(n1166), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[30]), .QN(n1165));
   SDFFARX1 \key_reg_reg[7][29]  (.D(n787), .SI(n1167), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[29]), .QN(n1166));
   SDFFARX1 \key_reg_reg[7][28]  (.D(n786), .SI(n1168), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[28]), .QN(n1167));
   SDFFARX1 \key_reg_reg[7][27]  (.D(n785), .SI(n1169), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[27]), .QN(n1168));
   SDFFARX1 \key_reg_reg[7][26]  (.D(n784), .SI(n1170), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[26]), .QN(n1169));
   SDFFARX1 \key_reg_reg[7][25]  (.D(n783), .SI(n1171), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[25]), .QN(n1170));
   SDFFARX1 \key_reg_reg[7][24]  (.D(n782), .SI(n1172), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[24]), .QN(n1171));
   SDFFARX1 \key_reg_reg[7][23]  (.D(n781), .SI(n1173), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[23]), .QN(n1172));
   SDFFARX1 \key_reg_reg[7][22]  (.D(n780), .SI(n1174), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1085), .Q(core_key[22]), .QN(n1173));
   SDFFARX1 \key_reg_reg[7][21]  (.D(n779), .SI(n1175), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[21]), .QN(n1174));
   SDFFARX1 \key_reg_reg[7][20]  (.D(n778), .SI(n1176), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[20]), .QN(n1175));
   SDFFARX1 \key_reg_reg[7][19]  (.D(n777), .SI(n1177), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[19]), .QN(n1176));
   SDFFARX1 \key_reg_reg[7][18]  (.D(n776), .SI(n1178), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[18]), .QN(n1177));
   SDFFARX1 \key_reg_reg[7][17]  (.D(n775), .SI(n1179), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[17]), .QN(n1178));
   SDFFARX1 \key_reg_reg[7][16]  (.D(n774), .SI(n1180), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[16]), .QN(n1179));
   SDFFARX1 \key_reg_reg[7][15]  (.D(n773), .SI(n1181), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[15]), .QN(n1180));
   SDFFARX1 \key_reg_reg[7][14]  (.D(n772), .SI(n1182), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[14]), .QN(n1181));
   SDFFARX1 \key_reg_reg[7][13]  (.D(n771), .SI(n1183), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[13]), .QN(n1182));
   SDFFARX1 \key_reg_reg[7][12]  (.D(n770), .SI(n1184), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[12]), .QN(n1183));
   SDFFARX1 \key_reg_reg[7][11]  (.D(n769), .SI(n1185), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[11]), .QN(n1184));
   SDFFARX1 \key_reg_reg[7][10]  (.D(n768), .SI(n1186), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1084), .Q(core_key[10]), .QN(n1185));
   SDFFARX1 \key_reg_reg[7][9]  (.D(n767), .SI(n1187), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[9]), .QN(n1186));
   SDFFARX1 \key_reg_reg[7][8]  (.D(n766), .SI(n1188), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[8]), .QN(n1187));
   SDFFARX1 \key_reg_reg[7][7]  (.D(n765), .SI(n1189), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[7]), .QN(n1188));
   SDFFARX1 \key_reg_reg[7][6]  (.D(n764), .SI(n1190), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[6]), .QN(n1189));
   SDFFARX1 \key_reg_reg[7][5]  (.D(n763), .SI(n1191), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[5]), .QN(n1190));
   SDFFARX1 \key_reg_reg[7][4]  (.D(n762), .SI(n1192), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[4]), .QN(n1191));
   SDFFARX1 \key_reg_reg[7][3]  (.D(n761), .SI(n1193), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[3]), .QN(n1192));
   SDFFARX1 \key_reg_reg[7][2]  (.D(n760), .SI(n1194), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[2]), .QN(n1193));
   SDFFARX1 \key_reg_reg[7][1]  (.D(n759), .SI(n1195), .SE(TEST_SE), .CLK(n1562), .RSTB(
          n1083), .Q(core_key[1]), .QN(n1194));
   SDFFARX1 \key_reg_reg[7][0]  (.D(n758), .SI(n1196), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1083), .Q(core_key[0]), .QN(n1195));
   SDFFARX1 next_reg_reg (.D(next_new), .SI(n1163), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1083), .Q(core_next), .QN(n1162));
   SDFFARX1 init_reg_reg (.D(init_new), .SI(n1421), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1083), .Q(core_init), .QN(n1420));
   SDFFARX1 keylen_reg_reg (.D(n757), .SI(n1164), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_keylen), .QN(n1163));
   SDFFARX1 encdec_reg_reg (.D(n756), .SI(n1422), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_encdec), .QN(n1421));
   SDFFARX1 \block_reg_reg[0][31]  (.D(n755), .SI(n1526), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[127]), .QN(n1525));
   SDFFARX1 \block_reg_reg[0][30]  (.D(n754), .SI(n1527), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[126]), .QN(n1526));
   SDFFARX1 \block_reg_reg[0][29]  (.D(n753), .SI(n1528), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[125]), .QN(n1527));
   SDFFARX1 \block_reg_reg[0][28]  (.D(n752), .SI(n1529), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[124]), .QN(n1528));
   SDFFARX1 \block_reg_reg[0][27]  (.D(n751), .SI(n1530), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[123]), .QN(n1529));
   SDFFARX1 \block_reg_reg[0][26]  (.D(n750), .SI(n1531), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[122]), .QN(n1530));
   SDFFARX1 \block_reg_reg[0][25]  (.D(n749), .SI(n1532), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[121]), .QN(n1531));
   SDFFARX1 \block_reg_reg[0][24]  (.D(n748), .SI(n1533), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[120]), .QN(n1532));
   SDFFARX1 \block_reg_reg[0][23]  (.D(n747), .SI(n1534), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[119]), .QN(n1533));
   SDFFARX1 \block_reg_reg[0][22]  (.D(n746), .SI(n1535), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1082), .Q(core_block[118]), .QN(n1534));
   SDFFARX1 \block_reg_reg[0][21]  (.D(n745), .SI(n1536), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[117]), .QN(n1535));
   SDFFARX1 \block_reg_reg[0][20]  (.D(n744), .SI(n1537), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[116]), .QN(n1536));
   SDFFARX1 \block_reg_reg[0][19]  (.D(n743), .SI(n1538), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[115]), .QN(n1537));
   SDFFARX1 \block_reg_reg[0][18]  (.D(n742), .SI(n1539), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[114]), .QN(n1538));
   SDFFARX1 \block_reg_reg[0][17]  (.D(n741), .SI(n1540), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[113]), .QN(n1539));
   SDFFARX1 \block_reg_reg[0][16]  (.D(n740), .SI(n1541), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[112]), .QN(n1540));
   SDFFARX1 \block_reg_reg[0][15]  (.D(n739), .SI(n1542), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[111]), .QN(n1541));
   SDFFARX1 \block_reg_reg[0][14]  (.D(n738), .SI(n1543), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[110]), .QN(n1542));
   SDFFARX1 \block_reg_reg[0][13]  (.D(n737), .SI(n1544), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[109]), .QN(n1543));
   SDFFARX1 \block_reg_reg[0][12]  (.D(n736), .SI(n1545), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[108]), .QN(n1544));
   SDFFARX1 \block_reg_reg[0][11]  (.D(n735), .SI(n1546), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[107]), .QN(n1545));
   SDFFARX1 \block_reg_reg[0][10]  (.D(n734), .SI(n1547), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1081), .Q(core_block[106]), .QN(n1546));
   SDFFARX1 \block_reg_reg[0][9]  (.D(n733), .SI(n1548), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[105]), .QN(n1547));
   SDFFARX1 \block_reg_reg[0][8]  (.D(n732), .SI(n1549), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[104]), .QN(n1548));
   SDFFARX1 \block_reg_reg[0][7]  (.D(n731), .SI(n1550), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[103]), .QN(n1549));
   SDFFARX1 \block_reg_reg[0][6]  (.D(n730), .SI(n1551), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[102]), .QN(n1550));
   SDFFARX1 \block_reg_reg[0][5]  (.D(n729), .SI(n1552), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[101]), .QN(n1551));
   SDFFARX1 \block_reg_reg[0][4]  (.D(n728), .SI(n1553), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[100]), .QN(n1552));
   SDFFARX1 \block_reg_reg[0][3]  (.D(n727), .SI(n1554), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[99]), .QN(n1553));
   SDFFARX1 \block_reg_reg[0][2]  (.D(n726), .SI(n1555), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[98]), .QN(n1554));
   SDFFARX1 \block_reg_reg[0][1]  (.D(n725), .SI(n1556), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[97]), .QN(n1555));
   SDFFARX1 \block_reg_reg[0][0]  (.D(n724), .SI(TEST_SI1), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[96]), .QN(n1556));
   SDFFARX1 \block_reg_reg[1][31]  (.D(n723), .SI(n1494), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[95]), .QN(n1493));
   SDFFARX1 \block_reg_reg[1][30]  (.D(n722), .SI(n1495), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1080), .Q(core_block[94]), .QN(n1494));
   SDFFARX1 \block_reg_reg[1][29]  (.D(n721), .SI(n1496), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[93]), .QN(n1495));
   SDFFARX1 \block_reg_reg[1][28]  (.D(n720), .SI(n1497), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[92]), .QN(n1496));
   SDFFARX1 \block_reg_reg[1][27]  (.D(n719), .SI(n1498), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[91]), .QN(n1497));
   SDFFARX1 \block_reg_reg[1][26]  (.D(n718), .SI(n1499), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[90]), .QN(n1498));
   SDFFARX1 \block_reg_reg[1][25]  (.D(n717), .SI(n1500), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[89]), .QN(n1499));
   SDFFARX1 \block_reg_reg[1][24]  (.D(n716), .SI(n1501), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[88]), .QN(n1500));
   SDFFARX1 \block_reg_reg[1][23]  (.D(n715), .SI(n1502), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[87]), .QN(n1501));
   SDFFARX1 \block_reg_reg[1][22]  (.D(n714), .SI(n1503), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[86]), .QN(n1502));
   SDFFARX1 \block_reg_reg[1][21]  (.D(n713), .SI(n1504), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[85]), .QN(n1503));
   SDFFARX1 \block_reg_reg[1][20]  (.D(n712), .SI(n1505), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[84]), .QN(n1504));
   SDFFARX1 \block_reg_reg[1][19]  (.D(n711), .SI(n1506), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[83]), .QN(n1505));
   SDFFARX1 \block_reg_reg[1][18]  (.D(n710), .SI(n1507), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1079), .Q(core_block[82]), .QN(n1506));
   SDFFARX1 \block_reg_reg[1][17]  (.D(n709), .SI(n1508), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1146), .Q(core_block[81]), .QN(n1507));
   SDFFARX1 \block_reg_reg[1][16]  (.D(n708), .SI(n1509), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[80]), .QN(n1508));
   SDFFARX1 \block_reg_reg[1][15]  (.D(n707), .SI(n1510), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[79]), .QN(n1509));
   SDFFARX1 \block_reg_reg[1][14]  (.D(n706), .SI(n1511), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[78]), .QN(n1510));
   SDFFARX1 \block_reg_reg[1][13]  (.D(n705), .SI(n1512), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[77]), .QN(n1511));
   SDFFARX1 \block_reg_reg[1][12]  (.D(n704), .SI(n1513), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[76]), .QN(n1512));
   SDFFARX1 \block_reg_reg[1][11]  (.D(n703), .SI(n1514), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[75]), .QN(n1513));
   SDFFARX1 \block_reg_reg[1][10]  (.D(n702), .SI(n1515), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[74]), .QN(n1514));
   SDFFARX1 \block_reg_reg[1][9]  (.D(n701), .SI(n1516), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[73]), .QN(n1515));
   SDFFARX1 \block_reg_reg[1][8]  (.D(n700), .SI(n1517), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[72]), .QN(n1516));
   SDFFARX1 \block_reg_reg[1][7]  (.D(n699), .SI(n1518), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[71]), .QN(n1517));
   SDFFARX1 \block_reg_reg[1][6]  (.D(n698), .SI(n1519), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[70]), .QN(n1518));
   SDFFARX1 \block_reg_reg[1][5]  (.D(n697), .SI(n1520), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1074), .Q(core_block[69]), .QN(n1519));
   SDFFARX1 \block_reg_reg[1][4]  (.D(n696), .SI(n1521), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[68]), .QN(n1520));
   SDFFARX1 \block_reg_reg[1][3]  (.D(n695), .SI(n1522), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[67]), .QN(n1521));
   SDFFARX1 \block_reg_reg[1][2]  (.D(n694), .SI(n1523), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[66]), .QN(n1522));
   SDFFARX1 \block_reg_reg[1][1]  (.D(n693), .SI(n1524), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[65]), .QN(n1523));
   SDFFARX1 \block_reg_reg[1][0]  (.D(n692), .SI(n1525), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[64]), .QN(n1524));
   SDFFARX1 \block_reg_reg[2][31]  (.D(n691), .SI(n1462), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[63]), .QN(n1461));
   SDFFARX1 \block_reg_reg[2][30]  (.D(n690), .SI(n1463), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[62]), .QN(n1462));
   SDFFARX1 \block_reg_reg[2][29]  (.D(n689), .SI(n1464), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[61]), .QN(n1463));
   SDFFARX1 \block_reg_reg[2][28]  (.D(n688), .SI(n1465), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[60]), .QN(n1464));
   SDFFARX1 \block_reg_reg[2][27]  (.D(n687), .SI(n1466), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[59]), .QN(n1465));
   SDFFARX1 \block_reg_reg[2][26]  (.D(n686), .SI(n1467), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[58]), .QN(n1466));
   SDFFARX1 \block_reg_reg[2][25]  (.D(n685), .SI(n1468), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1073), .Q(core_block[57]), .QN(n1467));
   SDFFARX1 \block_reg_reg[2][24]  (.D(n684), .SI(n1469), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[56]), .QN(n1468));
   SDFFARX1 \block_reg_reg[2][23]  (.D(n683), .SI(n1470), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[55]), .QN(n1469));
   SDFFARX1 \block_reg_reg[2][22]  (.D(n682), .SI(n1471), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[54]), .QN(n1470));
   SDFFARX1 \block_reg_reg[2][21]  (.D(n681), .SI(n1472), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[53]), .QN(n1471));
   SDFFARX1 \block_reg_reg[2][20]  (.D(n680), .SI(n1473), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[52]), .QN(n1472));
   SDFFARX1 \block_reg_reg[2][19]  (.D(n679), .SI(n1474), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[51]), .QN(n1473));
   SDFFARX1 \block_reg_reg[2][18]  (.D(n678), .SI(n1475), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[50]), .QN(n1474));
   SDFFARX1 \block_reg_reg[2][17]  (.D(n677), .SI(n1476), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[49]), .QN(n1475));
   SDFFARX1 \block_reg_reg[2][16]  (.D(n676), .SI(n1477), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[48]), .QN(n1476));
   SDFFARX1 \block_reg_reg[2][15]  (.D(n675), .SI(n1478), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[47]), .QN(n1477));
   SDFFARX1 \block_reg_reg[2][14]  (.D(n674), .SI(n1479), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[46]), .QN(n1478));
   SDFFARX1 \block_reg_reg[2][13]  (.D(n673), .SI(n1480), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1072), .Q(core_block[45]), .QN(n1479));
   SDFFARX1 \block_reg_reg[2][12]  (.D(n672), .SI(n1481), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[44]), .QN(n1480));
   SDFFARX1 \block_reg_reg[2][11]  (.D(n671), .SI(n1482), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[43]), .QN(n1481));
   SDFFARX1 \block_reg_reg[2][10]  (.D(n670), .SI(n1483), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[42]), .QN(n1482));
   SDFFARX1 \block_reg_reg[2][9]  (.D(n669), .SI(n1484), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[41]), .QN(n1483));
   SDFFARX1 \block_reg_reg[2][8]  (.D(n668), .SI(n1485), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[40]), .QN(n1484));
   SDFFARX1 \block_reg_reg[2][7]  (.D(n667), .SI(n1486), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[39]), .QN(n1485));
   SDFFARX1 \block_reg_reg[2][6]  (.D(n666), .SI(n1487), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[38]), .QN(n1486));
   SDFFARX1 \block_reg_reg[2][5]  (.D(n665), .SI(n1488), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[37]), .QN(n1487));
   SDFFARX1 \block_reg_reg[2][4]  (.D(n664), .SI(n1489), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[36]), .QN(n1488));
   SDFFARX1 \block_reg_reg[2][3]  (.D(n663), .SI(n1490), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[35]), .QN(n1489));
   SDFFARX1 \block_reg_reg[2][2]  (.D(n662), .SI(n1491), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[34]), .QN(n1490));
   SDFFARX1 \block_reg_reg[2][1]  (.D(n661), .SI(n1492), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1071), .Q(core_block[33]), .QN(n1491));
   SDFFARX1 \block_reg_reg[2][0]  (.D(n660), .SI(n1493), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[32]), .QN(n1492));
   SDFFARX1 \block_reg_reg[3][31]  (.D(n659), .SI(n1430), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[31]), .QN(n1429));
   SDFFARX1 \block_reg_reg[3][30]  (.D(n658), .SI(n1431), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[30]), .QN(n1430));
   SDFFARX1 \block_reg_reg[3][29]  (.D(n657), .SI(n1432), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[29]), .QN(n1431));
   SDFFARX1 \block_reg_reg[3][28]  (.D(n656), .SI(n1433), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[28]), .QN(n1432));
   SDFFARX1 \block_reg_reg[3][27]  (.D(n655), .SI(n1434), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[27]), .QN(n1433));
   SDFFARX1 \block_reg_reg[3][26]  (.D(n654), .SI(n1435), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[26]), .QN(n1434));
   SDFFARX1 \block_reg_reg[3][25]  (.D(n653), .SI(n1436), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[25]), .QN(n1435));
   SDFFARX1 \block_reg_reg[3][24]  (.D(n652), .SI(n1437), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[24]), .QN(n1436));
   SDFFARX1 \block_reg_reg[3][23]  (.D(n651), .SI(n1438), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[23]), .QN(n1437));
   SDFFARX1 \block_reg_reg[3][22]  (.D(n650), .SI(n1439), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[22]), .QN(n1438));
   SDFFARX1 \block_reg_reg[3][21]  (.D(n649), .SI(n1440), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1070), .Q(core_block[21]), .QN(n1439));
   SDFFARX1 \block_reg_reg[3][20]  (.D(n648), .SI(n1441), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[20]), .QN(n1440));
   SDFFARX1 \block_reg_reg[3][19]  (.D(n647), .SI(n1442), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[19]), .QN(n1441));
   SDFFARX1 \block_reg_reg[3][18]  (.D(n646), .SI(n1443), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[18]), .QN(n1442));
   SDFFARX1 \block_reg_reg[3][17]  (.D(n645), .SI(n1444), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[17]), .QN(n1443));
   SDFFARX1 \block_reg_reg[3][16]  (.D(n644), .SI(n1445), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[16]), .QN(n1444));
   SDFFARX1 \block_reg_reg[3][15]  (.D(n643), .SI(n1446), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[15]), .QN(n1445));
   SDFFARX1 \block_reg_reg[3][14]  (.D(n642), .SI(n1447), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[14]), .QN(n1446));
   SDFFARX1 \block_reg_reg[3][13]  (.D(n641), .SI(n1448), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[13]), .QN(n1447));
   SDFFARX1 \block_reg_reg[3][12]  (.D(n640), .SI(n1449), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[12]), .QN(n1448));
   SDFFARX1 \block_reg_reg[3][11]  (.D(n639), .SI(n1450), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[11]), .QN(n1449));
   SDFFARX1 \block_reg_reg[3][10]  (.D(n638), .SI(n1451), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[10]), .QN(n1450));
   SDFFARX1 \block_reg_reg[3][9]  (.D(n637), .SI(n1452), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1069), .Q(core_block[9]), .QN(n1451));
   SDFFARX1 \block_reg_reg[3][8]  (.D(n636), .SI(n1453), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[8]), .QN(n1452));
   SDFFARX1 \block_reg_reg[3][7]  (.D(n635), .SI(n1454), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[7]), .QN(n1453));
   SDFFARX1 \block_reg_reg[3][6]  (.D(n634), .SI(n1455), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[6]), .QN(n1454));
   SDFFARX1 \block_reg_reg[3][5]  (.D(n633), .SI(n1456), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[5]), .QN(n1455));
   SDFFARX1 \block_reg_reg[3][4]  (.D(n632), .SI(n1457), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[4]), .QN(n1456));
   SDFFARX1 \block_reg_reg[3][3]  (.D(n631), .SI(n1458), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[3]), .QN(n1457));
   SDFFARX1 \block_reg_reg[3][2]  (.D(n630), .SI(n1459), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[2]), .QN(n1458));
   SDFFARX1 \block_reg_reg[3][1]  (.D(n629), .SI(n1460), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[1]), .QN(n1459));
   SDFFARX1 \block_reg_reg[3][0]  (.D(n628), .SI(n1461), .SE(TEST_SE_buf_net0), .CLK(
          n1562_buf_net0), .RSTB(n1068), .Q(core_block[0]), .QN(n1460));
   SDFFARX1 valid_reg_reg (.D(core_valid), .SI(result_reg[127]), .SE(TEST_SE_buf_net0), .
          CLK(n1562_buf_net0), .RSTB(n1068), .Q(valid_reg));
   SDFFARX1 \result_reg_reg[0]  (.D(core_result[0]), .SI(ready_reg), .SE(TEST_SE_buf_net0)
          , .CLK(n1562_buf_net0), .RSTB(n1068), .Q(result_reg[0]));
   SDFFARX1 \result_reg_reg[1]  (.D(core_result[1]), .SI(result_reg[0]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1068), .Q(result_reg[1]));
   SDFFARX1 \result_reg_reg[2]  (.D(core_result[2]), .SI(result_reg[1]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[2]));
   SDFFARX1 \result_reg_reg[3]  (.D(core_result[3]), .SI(result_reg[2]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[3]));
   SDFFARX1 \result_reg_reg[4]  (.D(core_result[4]), .SI(result_reg[3]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[4]));
   SDFFARX1 \result_reg_reg[5]  (.D(core_result[5]), .SI(result_reg[4]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[5]));
   SDFFARX1 \result_reg_reg[6]  (.D(core_result[6]), .SI(result_reg[5]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[6]));
   SDFFARX1 \result_reg_reg[7]  (.D(core_result[7]), .SI(result_reg[6]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[7]));
   SDFFARX1 \result_reg_reg[8]  (.D(core_result[8]), .SI(result_reg[7]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[8]));
   SDFFARX1 \result_reg_reg[9]  (.D(core_result[9]), .SI(result_reg[8]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[9]));
   SDFFARX1 \result_reg_reg[10]  (.D(core_result[10]), .SI(result_reg[9]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[10]));
   SDFFARX1 \result_reg_reg[11]  (.D(core_result[11]), .SI(result_reg[10]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[11]));
   SDFFARX1 \result_reg_reg[12]  (.D(core_result[12]), .SI(result_reg[11]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[12]));
   SDFFARX1 \result_reg_reg[13]  (.D(core_result[13]), .SI(result_reg[12]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1067), .Q(result_reg[13]));
   SDFFARX1 \result_reg_reg[14]  (.D(core_result[14]), .SI(result_reg[13]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[14]));
   SDFFARX1 \result_reg_reg[15]  (.D(core_result[15]), .SI(result_reg[14]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[15]));
   SDFFARX1 \result_reg_reg[16]  (.D(core_result[16]), .SI(result_reg[15]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[16]));
   SDFFARX1 \result_reg_reg[17]  (.D(core_result[17]), .SI(result_reg[16]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[17]));
   SDFFARX1 \result_reg_reg[18]  (.D(core_result[18]), .SI(result_reg[17]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[18]));
   SDFFARX1 \result_reg_reg[19]  (.D(core_result[19]), .SI(result_reg[18]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[19]));
   SDFFARX1 \result_reg_reg[20]  (.D(core_result[20]), .SI(result_reg[19]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[20]));
   SDFFARX1 \result_reg_reg[21]  (.D(core_result[21]), .SI(result_reg[20]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[21]));
   SDFFARX1 \result_reg_reg[22]  (.D(core_result[22]), .SI(result_reg[21]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[22]));
   SDFFARX1 \result_reg_reg[23]  (.D(core_result[23]), .SI(result_reg[22]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[23]));
   SDFFARX1 \result_reg_reg[24]  (.D(core_result[24]), .SI(result_reg[23]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[24]));
   SDFFARX1 \result_reg_reg[25]  (.D(core_result[25]), .SI(result_reg[24]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1066), .Q(result_reg[25]));
   SDFFARX1 \result_reg_reg[26]  (.D(core_result[26]), .SI(result_reg[25]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[26]));
   SDFFARX1 \result_reg_reg[27]  (.D(core_result[27]), .SI(result_reg[26]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[27]));
   SDFFARX1 \result_reg_reg[28]  (.D(core_result[28]), .SI(result_reg[27]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[28]));
   SDFFARX1 \result_reg_reg[29]  (.D(core_result[29]), .SI(result_reg[28]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[29]));
   SDFFARX1 \result_reg_reg[30]  (.D(core_result[30]), .SI(result_reg[29]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[30]));
   SDFFARX1 \result_reg_reg[31]  (.D(core_result[31]), .SI(result_reg[30]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[31]));
   SDFFARX1 \result_reg_reg[32]  (.D(core_result[32]), .SI(result_reg[31]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[32]));
   SDFFARX1 \result_reg_reg[33]  (.D(core_result[33]), .SI(result_reg[32]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[33]));
   SDFFARX1 \result_reg_reg[34]  (.D(core_result[34]), .SI(result_reg[33]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[34]));
   SDFFARX1 \result_reg_reg[35]  (.D(core_result[35]), .SI(result_reg[34]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[35]));
   SDFFARX1 \result_reg_reg[36]  (.D(core_result[36]), .SI(result_reg[35]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[36]));
   SDFFARX1 \result_reg_reg[37]  (.D(core_result[37]), .SI(result_reg[36]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1065), .Q(result_reg[37]));
   SDFFARX1 \result_reg_reg[38]  (.D(core_result[38]), .SI(result_reg[37]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[38]));
   SDFFARX1 \result_reg_reg[39]  (.D(core_result[39]), .SI(result_reg[38]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[39]));
   SDFFARX1 \result_reg_reg[40]  (.D(core_result[40]), .SI(result_reg[39]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[40]));
   SDFFARX1 \result_reg_reg[41]  (.D(core_result[41]), .SI(result_reg[40]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[41]));
   SDFFARX1 \result_reg_reg[42]  (.D(core_result[42]), .SI(result_reg[41]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[42]));
   SDFFARX1 \result_reg_reg[43]  (.D(core_result[43]), .SI(result_reg[42]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[43]));
   SDFFARX1 \result_reg_reg[44]  (.D(core_result[44]), .SI(result_reg[43]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[44]));
   SDFFARX1 \result_reg_reg[45]  (.D(core_result[45]), .SI(result_reg[44]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[45]));
   SDFFARX1 \result_reg_reg[46]  (.D(core_result[46]), .SI(result_reg[45]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[46]));
   SDFFARX1 \result_reg_reg[47]  (.D(core_result[47]), .SI(result_reg[46]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[47]));
   SDFFARX1 \result_reg_reg[48]  (.D(core_result[48]), .SI(result_reg[47]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[48]));
   SDFFARX1 \result_reg_reg[49]  (.D(core_result[49]), .SI(result_reg[48]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1018), .Q(result_reg[49]));
   SDFFARX1 \result_reg_reg[50]  (.D(core_result[50]), .SI(result_reg[49]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[50]));
   SDFFARX1 \result_reg_reg[51]  (.D(core_result[51]), .SI(result_reg[50]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[51]));
   SDFFARX1 \result_reg_reg[52]  (.D(core_result[52]), .SI(result_reg[51]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[52]));
   SDFFARX1 \result_reg_reg[53]  (.D(core_result[53]), .SI(result_reg[52]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[53]));
   SDFFARX1 \result_reg_reg[54]  (.D(core_result[54]), .SI(result_reg[53]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[54]));
   SDFFARX1 \result_reg_reg[55]  (.D(core_result[55]), .SI(result_reg[54]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[55]));
   SDFFARX1 \result_reg_reg[56]  (.D(core_result[56]), .SI(result_reg[55]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[56]));
   SDFFARX1 \result_reg_reg[57]  (.D(core_result[57]), .SI(result_reg[56]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[57]));
   SDFFARX1 \result_reg_reg[58]  (.D(core_result[58]), .SI(result_reg[57]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[58]));
   SDFFARX1 \result_reg_reg[59]  (.D(core_result[59]), .SI(result_reg[58]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[59]));
   SDFFARX1 \result_reg_reg[60]  (.D(core_result[60]), .SI(result_reg[59]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[60]));
   SDFFARX1 \result_reg_reg[61]  (.D(core_result[61]), .SI(result_reg[60]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1019), .Q(result_reg[61]));
   SDFFARX1 \result_reg_reg[62]  (.D(core_result[62]), .SI(result_reg[61]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[62]));
   SDFFARX1 \result_reg_reg[63]  (.D(core_result[63]), .SI(result_reg[62]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[63]));
   SDFFARX1 \result_reg_reg[64]  (.D(core_result[64]), .SI(result_reg[63]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[64]));
   SDFFARX1 \result_reg_reg[65]  (.D(core_result[65]), .SI(result_reg[64]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[65]));
   SDFFARX1 \result_reg_reg[66]  (.D(core_result[66]), .SI(result_reg[65]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[66]));
   SDFFARX1 \result_reg_reg[67]  (.D(core_result[67]), .SI(result_reg[66]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[67]));
   SDFFARX1 \result_reg_reg[68]  (.D(core_result[68]), .SI(result_reg[67]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[68]));
   SDFFARX1 \result_reg_reg[69]  (.D(core_result[69]), .SI(result_reg[68]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[69]));
   SDFFARX1 \result_reg_reg[70]  (.D(core_result[70]), .SI(result_reg[69]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[70]));
   SDFFARX1 \result_reg_reg[71]  (.D(core_result[71]), .SI(result_reg[70]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[71]));
   SDFFARX1 \result_reg_reg[72]  (.D(core_result[72]), .SI(result_reg[71]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[72]));
   SDFFARX1 \result_reg_reg[73]  (.D(core_result[73]), .SI(result_reg[72]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1020), .Q(result_reg[73]));
   SDFFARX1 \result_reg_reg[74]  (.D(core_result[74]), .SI(result_reg[73]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[74]));
   SDFFARX1 \result_reg_reg[75]  (.D(core_result[75]), .SI(result_reg[74]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[75]));
   SDFFARX1 \result_reg_reg[76]  (.D(core_result[76]), .SI(result_reg[75]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[76]));
   SDFFARX1 \result_reg_reg[77]  (.D(core_result[77]), .SI(result_reg[76]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[77]));
   SDFFARX1 \result_reg_reg[78]  (.D(core_result[78]), .SI(result_reg[77]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[78]));
   SDFFARX1 \result_reg_reg[79]  (.D(core_result[79]), .SI(result_reg[78]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[79]));
   SDFFARX1 \result_reg_reg[80]  (.D(core_result[80]), .SI(result_reg[79]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[80]));
   SDFFARX1 \result_reg_reg[81]  (.D(core_result[81]), .SI(result_reg[80]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[81]));
   SDFFARX1 \result_reg_reg[82]  (.D(core_result[82]), .SI(result_reg[81]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[82]));
   SDFFARX1 \result_reg_reg[83]  (.D(core_result[83]), .SI(result_reg[82]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[83]));
   SDFFARX1 \result_reg_reg[84]  (.D(core_result[84]), .SI(result_reg[83]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[84]));
   SDFFARX1 \result_reg_reg[85]  (.D(core_result[85]), .SI(result_reg[84]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1021), .Q(result_reg[85]));
   SDFFARX1 \result_reg_reg[86]  (.D(core_result[86]), .SI(result_reg[85]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[86]));
   SDFFARX1 \result_reg_reg[87]  (.D(core_result[87]), .SI(result_reg[86]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[87]));
   SDFFARX1 \result_reg_reg[88]  (.D(core_result[88]), .SI(result_reg[87]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[88]));
   SDFFARX1 \result_reg_reg[89]  (.D(core_result[89]), .SI(result_reg[88]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[89]));
   SDFFARX1 \result_reg_reg[90]  (.D(core_result[90]), .SI(result_reg[89]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[90]));
   SDFFARX1 \result_reg_reg[91]  (.D(core_result[91]), .SI(result_reg[90]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[91]));
   SDFFARX1 \result_reg_reg[92]  (.D(core_result[92]), .SI(result_reg[91]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[92]));
   SDFFARX1 \result_reg_reg[93]  (.D(core_result[93]), .SI(result_reg[92]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[93]));
   SDFFARX1 \result_reg_reg[94]  (.D(core_result[94]), .SI(result_reg[93]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[94]));
   SDFFARX1 \result_reg_reg[95]  (.D(core_result[95]), .SI(result_reg[94]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[95]));
   SDFFARX1 \result_reg_reg[96]  (.D(core_result[96]), .SI(result_reg[95]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[96]));
   SDFFARX1 \result_reg_reg[97]  (.D(core_result[97]), .SI(result_reg[96]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1022), .Q(result_reg[97]));
   SDFFARX1 \result_reg_reg[98]  (.D(core_result[98]), .SI(result_reg[97]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[98]));
   SDFFARX1 \result_reg_reg[99]  (.D(core_result[99]), .SI(result_reg[98]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[99]));
   SDFFARX1 \result_reg_reg[100]  (.D(core_result[100]), .SI(result_reg[99]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[100]));
   SDFFARX1 \result_reg_reg[101]  (.D(core_result[101]), .SI(result_reg[100]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[101]));
   SDFFARX1 \result_reg_reg[102]  (.D(core_result[102]), .SI(result_reg[101]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[102]));
   SDFFARX1 \result_reg_reg[103]  (.D(core_result[103]), .SI(result_reg[102]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[103]));
   SDFFARX1 \result_reg_reg[104]  (.D(core_result[104]), .SI(result_reg[103]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[104]));
   SDFFARX1 \result_reg_reg[105]  (.D(core_result[105]), .SI(result_reg[104]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[105]));
   SDFFARX1 \result_reg_reg[106]  (.D(core_result[106]), .SI(result_reg[105]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[106]));
   SDFFARX1 \result_reg_reg[107]  (.D(core_result[107]), .SI(result_reg[106]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[107]));
   SDFFARX1 \result_reg_reg[108]  (.D(core_result[108]), .SI(result_reg[107]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[108]));
   SDFFARX1 \result_reg_reg[109]  (.D(core_result[109]), .SI(result_reg[108]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1023), .Q(result_reg[109]));
   SDFFARX1 \result_reg_reg[110]  (.D(core_result[110]), .SI(result_reg[109]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[110]));
   SDFFARX1 \result_reg_reg[111]  (.D(core_result[111]), .SI(result_reg[110]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[111]));
   SDFFARX1 \result_reg_reg[112]  (.D(core_result[112]), .SI(result_reg[111]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[112]));
   SDFFARX1 \result_reg_reg[113]  (.D(core_result[113]), .SI(result_reg[112]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[113]));
   SDFFARX1 \result_reg_reg[114]  (.D(core_result[114]), .SI(result_reg[113]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[114]));
   SDFFARX1 \result_reg_reg[115]  (.D(core_result[115]), .SI(result_reg[114]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[115]));
   SDFFARX1 \result_reg_reg[116]  (.D(core_result[116]), .SI(result_reg[115]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[116]));
   SDFFARX1 \result_reg_reg[117]  (.D(core_result[117]), .SI(result_reg[116]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[117]));
   SDFFARX1 \result_reg_reg[118]  (.D(core_result[118]), .SI(result_reg[117]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[118]));
   SDFFARX1 \result_reg_reg[119]  (.D(core_result[119]), .SI(result_reg[118]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[119]));
   SDFFARX1 \result_reg_reg[120]  (.D(core_result[120]), .SI(result_reg[119]), .SE(
          TEST_SE_buf_net0), .CLK(n1562_buf_net0), .RSTB(n1024), .Q(result_reg[120]));
   SDFFARX1 \result_reg_reg[121]  (.D(core_result[121]), .SI(result_reg[120]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1024), .Q(result_reg[121]));
   SDFFARX1 \result_reg_reg[122]  (.D(core_result[122]), .SI(result_reg[121]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[122]));
   SDFFARX1 \result_reg_reg[123]  (.D(core_result[123]), .SI(result_reg[122]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[123]));
   SDFFARX1 \result_reg_reg[124]  (.D(core_result[124]), .SI(result_reg[123]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[124]));
   SDFFARX1 \result_reg_reg[125]  (.D(core_result[125]), .SI(result_reg[124]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[125]));
   SDFFARX1 \result_reg_reg[126]  (.D(core_result[126]), .SI(result_reg[125]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[126]));
   SDFFARX1 \result_reg_reg[127]  (.D(core_result[127]), .SI(result_reg[126]), .SE(
          TEST_SE_buf_net1), .CLK(n1562_buf_net1), .RSTB(n1025), .Q(result_reg[127]));
   SDFFARX1 ready_reg_reg (.D(core_ready), .SI(n1162), .SE(TEST_SE_buf_net1), .CLK(
          n1562_buf_net1), .RSTB(n1025), .Q(ready_reg));
   AO221X1 U570 (.IN1(result_reg[73]), .IN2(n1140), .IN3(result_reg[105]), .IN4(n1137), .
          IN5(n552), .Q(read_data[9]));
   AO221X1 U571 (.IN1(result_reg[9]), .IN2(n1134), .IN3(result_reg[41]), .IN4(n1131), .IN5(
          n555), .Q(n552));
   AO221X1 U572 (.IN1(result_reg[72]), .IN2(n1142), .IN3(result_reg[104]), .IN4(n1138), .
          IN5(n556), .Q(read_data[8]));
   AO221X1 U573 (.IN1(result_reg[8]), .IN2(n1136), .IN3(result_reg[40]), .IN4(n1133), .IN5(
          n557), .Q(n556));
   AO221X1 U574 (.IN1(result_reg[7]), .IN2(n1136), .IN3(result_reg[39]), .IN4(n1133), .IN5(
          n558), .Q(read_data[7]));
   AO22X1 U575 (.IN1(result_reg[103]), .IN2(n1139), .IN3(result_reg[71]), .IN4(n1140), .Q(
          n558));
   AO221X1 U576 (.IN1(result_reg[6]), .IN2(n1136), .IN3(result_reg[38]), .IN4(n1133), .IN5(
          n559), .Q(read_data[6]));
   AO22X1 U577 (.IN1(result_reg[102]), .IN2(n1139), .IN3(result_reg[70]), .IN4(n1140), .Q(
          n559));
   AO221X1 U578 (.IN1(result_reg[69]), .IN2(n1142), .IN3(result_reg[101]), .IN4(n1138), .
          IN5(n560), .Q(read_data[5]));
   AO221X1 U579 (.IN1(result_reg[5]), .IN2(n1135), .IN3(result_reg[37]), .IN4(n1132), .IN5(
          n561), .Q(n560));
   AO221X1 U580 (.IN1(result_reg[68]), .IN2(n1142), .IN3(result_reg[100]), .IN4(n1138), .
          IN5(n562), .Q(read_data[4]));
   AO221X1 U581 (.IN1(result_reg[4]), .IN2(n1136), .IN3(result_reg[36]), .IN4(n1133), .IN5(
          n563), .Q(n562));
   AO221X1 U582 (.IN1(result_reg[67]), .IN2(n1142), .IN3(result_reg[99]), .IN4(n1138), .
          IN5(n564), .Q(read_data[3]));
   AO221X1 U584 (.IN1(result_reg[31]), .IN2(n1135), .IN3(result_reg[63]), .IN4(n1132), .
          IN5(n566), .Q(read_data[31]));
   AO22X1 U585 (.IN1(result_reg[127]), .IN2(n1139), .IN3(result_reg[95]), .IN4(n1140), .Q(
          n566));
   AO221X1 U586 (.IN1(result_reg[94]), .IN2(n1142), .IN3(result_reg[126]), .IN4(n1138), .
          IN5(n567), .Q(read_data[30]));
   AO221X1 U587 (.IN1(result_reg[30]), .IN2(n1135), .IN3(result_reg[62]), .IN4(n1132), .
          IN5(n557), .Q(n567));
   AO221X1 U588 (.IN1(result_reg[66]), .IN2(n1142), .IN3(result_reg[98]), .IN4(n1138), .
          IN5(n568), .Q(read_data[2]));
   AO221X1 U590 (.IN1(result_reg[93]), .IN2(n1141), .IN3(result_reg[125]), .IN4(n1138), .
          IN5(n569), .Q(read_data[29]));
   AO221X1 U591 (.IN1(result_reg[29]), .IN2(n1135), .IN3(result_reg[61]), .IN4(n1132), .
          IN5(n561), .Q(n569));
   AO221X1 U592 (.IN1(result_reg[92]), .IN2(n1141), .IN3(result_reg[124]), .IN4(n1138), .
          IN5(n570), .Q(read_data[28]));
   AO221X1 U593 (.IN1(result_reg[28]), .IN2(n1135), .IN3(result_reg[60]), .IN4(n1132), .
          IN5(n563), .Q(n570));
   AO221X1 U594 (.IN1(result_reg[27]), .IN2(n1135), .IN3(result_reg[59]), .IN4(n1132), .
          IN5(n571), .Q(read_data[27]));
   AO22X1 U595 (.IN1(result_reg[123]), .IN2(n1138), .IN3(result_reg[91]), .IN4(n1140), .Q(
          n571));
   AO221X1 U596 (.IN1(result_reg[26]), .IN2(n1135), .IN3(result_reg[58]), .IN4(n1132), .
          IN5(n572), .Q(read_data[26]));
   AO22X1 U597 (.IN1(result_reg[122]), .IN2(n1138), .IN3(result_reg[90]), .IN4(n1140), .Q(
          n572));
   AO221X1 U598 (.IN1(result_reg[25]), .IN2(n1135), .IN3(result_reg[57]), .IN4(n1132), .
          IN5(n573), .Q(read_data[25]));
   AO22X1 U599 (.IN1(result_reg[121]), .IN2(n1138), .IN3(result_reg[89]), .IN4(n1140), .Q(
          n573));
   AO221X1 U600 (.IN1(result_reg[88]), .IN2(n1141), .IN3(result_reg[120]), .IN4(n1137), .
          IN5(n574), .Q(read_data[24]));
   AO221X1 U601 (.IN1(result_reg[24]), .IN2(n1135), .IN3(result_reg[56]), .IN4(n1132), .
          IN5(n557), .Q(n574));
   AO221X1 U602 (.IN1(result_reg[23]), .IN2(n1135), .IN3(result_reg[55]), .IN4(n1132), .
          IN5(n575), .Q(read_data[23]));
   AO22X1 U603 (.IN1(result_reg[119]), .IN2(n1138), .IN3(result_reg[87]), .IN4(n1140), .Q(
          n575));
   AO221X1 U604 (.IN1(result_reg[86]), .IN2(n1141), .IN3(result_reg[118]), .IN4(n1137), .
          IN5(n576), .Q(read_data[22]));
   AO221X1 U605 (.IN1(result_reg[22]), .IN2(n1135), .IN3(result_reg[54]), .IN4(n1132), .
          IN5(n557), .Q(n576));
   AO221X1 U606 (.IN1(result_reg[85]), .IN2(n1141), .IN3(result_reg[117]), .IN4(n1137), .
          IN5(n577), .Q(read_data[21]));
   AO221X1 U607 (.IN1(result_reg[21]), .IN2(n1134), .IN3(result_reg[53]), .IN4(n1131), .
          IN5(n561), .Q(n577));
   AO221X1 U608 (.IN1(result_reg[20]), .IN2(n1134), .IN3(result_reg[52]), .IN4(n1131), .
          IN5(n578), .Q(read_data[20]));
   AO22X1 U609 (.IN1(result_reg[116]), .IN2(n1138), .IN3(result_reg[84]), .IN4(n1140), .Q(
          n578));
   AOI222X1 U610 (.IN1(result_reg[1]), .IN2(n1136), .IN3(core_next), .IN4(n565), .IN5(
          valid_reg), .IN6(n581), .QN(n580));
   AOI222X1 U611 (.IN1(result_reg[97]), .IN2(n1139), .IN3(result_reg[33]), .IN4(n1133), .
          IN5(result_reg[65]), .IN6(n1140), .QN(n579));
   AO221X1 U612 (.IN1(result_reg[83]), .IN2(n1141), .IN3(result_reg[115]), .IN4(n1137), .
          IN5(n582), .Q(read_data[19]));
   AO221X1 U613 (.IN1(result_reg[19]), .IN2(n1134), .IN3(result_reg[51]), .IN4(n1131), .
          IN5(n563), .Q(n582));
   AO221X1 U614 (.IN1(result_reg[82]), .IN2(n1141), .IN3(result_reg[114]), .IN4(n1137), .
          IN5(n583), .Q(read_data[18]));
   AO221X1 U615 (.IN1(result_reg[18]), .IN2(n1134), .IN3(result_reg[50]), .IN4(n1131), .
          IN5(n555), .Q(n583));
   AO221X1 U616 (.IN1(result_reg[81]), .IN2(n1141), .IN3(result_reg[113]), .IN4(n1137), .
          IN5(n584), .Q(read_data[17]));
   AO221X1 U617 (.IN1(result_reg[17]), .IN2(n1135), .IN3(result_reg[49]), .IN4(n1132), .
          IN5(n563), .Q(n584));
   AO221X1 U618 (.IN1(result_reg[80]), .IN2(n1141), .IN3(result_reg[112]), .IN4(n1137), .
          IN5(n585), .Q(read_data[16]));
   AO221X1 U619 (.IN1(result_reg[16]), .IN2(n1134), .IN3(result_reg[48]), .IN4(n1131), .
          IN5(n557), .Q(n585));
   AO221X1 U620 (.IN1(result_reg[15]), .IN2(n1134), .IN3(result_reg[47]), .IN4(n1131), .
          IN5(n586), .Q(read_data[15]));
   AO22X1 U621 (.IN1(result_reg[111]), .IN2(n1139), .IN3(result_reg[79]), .IN4(n1140), .Q(
          n586));
   AO221X1 U622 (.IN1(result_reg[78]), .IN2(n1141), .IN3(result_reg[110]), .IN4(n1137), .
          IN5(n587), .Q(read_data[14]));
   AO221X1 U623 (.IN1(result_reg[14]), .IN2(n1134), .IN3(result_reg[46]), .IN4(n1131), .
          IN5(n557), .Q(n587));
   NOR3X0 U624 (.IN1(n588), .IN2(address[1]), .IN3(n589), .QN(n557));
   AO221X1 U625 (.IN1(result_reg[77]), .IN2(n1141), .IN3(result_reg[109]), .IN4(n1137), .
          IN5(n590), .Q(read_data[13]));
   AO221X1 U626 (.IN1(result_reg[13]), .IN2(n1134), .IN3(result_reg[45]), .IN4(n1131), .
          IN5(n561), .Q(n590));
   AOI21X1 U627 (.IN1(n589), .IN2(n591), .IN3(n588), .QN(n561));
   NAND3X0 U628 (.IN1(n1160), .IN2(n1158), .IN3(n592), .QN(n591));
   AO221X1 U629 (.IN1(result_reg[76]), .IN2(n1141), .IN3(result_reg[108]), .IN4(n1137), .
          IN5(n593), .Q(read_data[12]));
   AO221X1 U630 (.IN1(result_reg[12]), .IN2(n1134), .IN3(result_reg[44]), .IN4(n1131), .
          IN5(n555), .Q(n593));
   AO221X1 U631 (.IN1(result_reg[11]), .IN2(n1134), .IN3(result_reg[43]), .IN4(n1131), .
          IN5(n594), .Q(read_data[11]));
   AO22X1 U632 (.IN1(result_reg[107]), .IN2(n1139), .IN3(result_reg[75]), .IN4(n1140), .Q(
          n594));
   AO221X1 U633 (.IN1(result_reg[74]), .IN2(n1141), .IN3(result_reg[106]), .IN4(n1137), .
          IN5(n595), .Q(read_data[10]));
   AO221X1 U634 (.IN1(result_reg[10]), .IN2(n1134), .IN3(result_reg[42]), .IN4(n1131), .
          IN5(n563), .Q(n595));
   NOR3X0 U635 (.IN1(n589), .IN2(n588), .IN3(n1160), .QN(n563));
   NAND3X0 U636 (.IN1(n1161), .IN2(n1158), .IN3(n592), .QN(n589));
   AOI222X1 U637 (.IN1(result_reg[0]), .IN2(n1136), .IN3(core_init), .IN4(n565), .IN5(
          ready_reg), .IN6(n581), .QN(n597));
   AND4X1 U638 (.IN1(address[3]), .IN2(n598), .IN3(n1155), .IN4(n592), .Q(n581));
   NAND3X0 U639 (.IN1(cs), .IN2(n600), .IN3(we), .QN(n588));
   AOI222X1 U641 (.IN1(result_reg[96]), .IN2(n1139), .IN3(result_reg[32]), .IN4(n1133), .
          IN5(result_reg[64]), .IN6(n1140), .QN(n596));
   NOR3X0 U645 (.IN1(n1156), .IN2(n1154), .IN3(n600), .QN(n602));
   AND3X1 U646 (.IN1(write_data[1]), .IN2(n1157), .IN3(n606), .Q(next_new));
   AO22X1 U647 (.IN1(write_data[0]), .IN2(n1062), .IN3(core_block[0]), .IN4(n607), .Q(n628)
          );
   AO22X1 U648 (.IN1(n1062), .IN2(write_data[1]), .IN3(core_block[1]), .IN4(n607), .Q(n629)
          );
   AO22X1 U649 (.IN1(write_data[2]), .IN2(n1064), .IN3(core_block[2]), .IN4(n607), .Q(n630)
          );
   AO22X1 U650 (.IN1(write_data[3]), .IN2(n1064), .IN3(core_block[3]), .IN4(n607), .Q(n631)
          );
   AO22X1 U651 (.IN1(write_data[4]), .IN2(n1064), .IN3(core_block[4]), .IN4(n607), .Q(n632)
          );
   AO22X1 U652 (.IN1(write_data[5]), .IN2(n1064), .IN3(core_block[5]), .IN4(n607), .Q(n633)
          );
   AO22X1 U653 (.IN1(write_data[6]), .IN2(n1064), .IN3(core_block[6]), .IN4(n607), .Q(n634)
          );
   AO22X1 U654 (.IN1(write_data[7]), .IN2(n1064), .IN3(core_block[7]), .IN4(n607), .Q(n635)
          );
   AO22X1 U655 (.IN1(write_data[8]), .IN2(n1064), .IN3(core_block[8]), .IN4(n1130), .Q(
          n636));
   AO22X1 U656 (.IN1(write_data[9]), .IN2(n1064), .IN3(core_block[9]), .IN4(n1130), .Q(
          n637));
   AO22X1 U657 (.IN1(write_data[10]), .IN2(n1063), .IN3(core_block[10]), .IN4(n1130), .Q(
          n638));
   AO22X1 U658 (.IN1(write_data[11]), .IN2(n1063), .IN3(core_block[11]), .IN4(n1130), .Q(
          n639));
   AO22X1 U659 (.IN1(write_data[12]), .IN2(n1063), .IN3(core_block[12]), .IN4(n1130), .Q(
          n640));
   AO22X1 U660 (.IN1(write_data[13]), .IN2(n1063), .IN3(core_block[13]), .IN4(n1130), .Q(
          n641));
   AO22X1 U661 (.IN1(write_data[14]), .IN2(n1063), .IN3(core_block[14]), .IN4(n1130), .Q(
          n642));
   AO22X1 U662 (.IN1(write_data[15]), .IN2(n1063), .IN3(core_block[15]), .IN4(n1130), .Q(
          n643));
   AO22X1 U663 (.IN1(write_data[16]), .IN2(n1063), .IN3(core_block[16]), .IN4(n1130), .Q(
          n644));
   AO22X1 U664 (.IN1(write_data[17]), .IN2(n1063), .IN3(core_block[17]), .IN4(n1130), .Q(
          n645));
   AO22X1 U665 (.IN1(write_data[18]), .IN2(n1063), .IN3(core_block[18]), .IN4(n1130), .Q(
          n646));
   AO22X1 U666 (.IN1(write_data[19]), .IN2(n1063), .IN3(core_block[19]), .IN4(n1130), .Q(
          n647));
   AO22X1 U667 (.IN1(write_data[20]), .IN2(n1063), .IN3(core_block[20]), .IN4(n1129), .Q(
          n648));
   AO22X1 U668 (.IN1(write_data[21]), .IN2(n1062), .IN3(core_block[21]), .IN4(n1129), .Q(
          n649));
   AO22X1 U669 (.IN1(write_data[22]), .IN2(n1062), .IN3(core_block[22]), .IN4(n1129), .Q(
          n650));
   AO22X1 U670 (.IN1(write_data[23]), .IN2(n1062), .IN3(core_block[23]), .IN4(n1129), .Q(
          n651));
   AO22X1 U671 (.IN1(write_data[24]), .IN2(n1062), .IN3(core_block[24]), .IN4(n1129), .Q(
          n652));
   AO22X1 U672 (.IN1(write_data[25]), .IN2(n1062), .IN3(core_block[25]), .IN4(n1129), .Q(
          n653));
   AO22X1 U673 (.IN1(write_data[26]), .IN2(n1062), .IN3(core_block[26]), .IN4(n1129), .Q(
          n654));
   AO22X1 U674 (.IN1(write_data[27]), .IN2(n1062), .IN3(core_block[27]), .IN4(n1129), .Q(
          n655));
   AO22X1 U675 (.IN1(write_data[28]), .IN2(n1062), .IN3(core_block[28]), .IN4(n1129), .Q(
          n656));
   AO22X1 U676 (.IN1(write_data[29]), .IN2(n1062), .IN3(core_block[29]), .IN4(n1129), .Q(
          n657));
   AO22X1 U677 (.IN1(write_data[30]), .IN2(n1062), .IN3(core_block[30]), .IN4(n1129), .Q(
          n658));
   AO22X1 U678 (.IN1(write_data[31]), .IN2(n1063), .IN3(core_block[31]), .IN4(n1129), .Q(
          n659));
   AO22X1 U679 (.IN1(n1059), .IN2(write_data[0]), .IN3(core_block[32]), .IN4(n610), .Q(
          n660));
   AO22X1 U680 (.IN1(n1059), .IN2(write_data[1]), .IN3(core_block[33]), .IN4(n610), .Q(
          n661));
   AO22X1 U681 (.IN1(n1059), .IN2(write_data[2]), .IN3(core_block[34]), .IN4(n610), .Q(
          n662));
   AO22X1 U682 (.IN1(n1059), .IN2(write_data[3]), .IN3(core_block[35]), .IN4(n610), .Q(
          n663));
   AO22X1 U683 (.IN1(n1059), .IN2(write_data[4]), .IN3(core_block[36]), .IN4(n610), .Q(
          n664));
   AO22X1 U684 (.IN1(n1059), .IN2(write_data[5]), .IN3(core_block[37]), .IN4(n610), .Q(
          n665));
   AO22X1 U685 (.IN1(n1059), .IN2(write_data[6]), .IN3(core_block[38]), .IN4(n610), .Q(
          n666));
   AO22X1 U686 (.IN1(n1059), .IN2(write_data[7]), .IN3(core_block[39]), .IN4(n610), .Q(
          n667));
   AO22X1 U687 (.IN1(n1059), .IN2(write_data[8]), .IN3(core_block[40]), .IN4(n1128), .Q(
          n668));
   AO22X1 U688 (.IN1(n1059), .IN2(write_data[9]), .IN3(core_block[41]), .IN4(n1128), .Q(
          n669));
   AO22X1 U689 (.IN1(n1059), .IN2(write_data[10]), .IN3(core_block[42]), .IN4(n1128), .Q(
          n670));
   AO22X1 U690 (.IN1(n1059), .IN2(write_data[11]), .IN3(core_block[43]), .IN4(n1128), .Q(
          n671));
   AO22X1 U691 (.IN1(n1060), .IN2(write_data[12]), .IN3(core_block[44]), .IN4(n1128), .Q(
          n672));
   AO22X1 U692 (.IN1(n1060), .IN2(write_data[13]), .IN3(core_block[45]), .IN4(n1128), .Q(
          n673));
   AO22X1 U693 (.IN1(n1060), .IN2(write_data[14]), .IN3(core_block[46]), .IN4(n1128), .Q(
          n674));
   AO22X1 U694 (.IN1(n1060), .IN2(write_data[15]), .IN3(core_block[47]), .IN4(n1128), .Q(
          n675));
   AO22X1 U695 (.IN1(n1060), .IN2(write_data[16]), .IN3(core_block[48]), .IN4(n1128), .Q(
          n676));
   AO22X1 U696 (.IN1(n1060), .IN2(write_data[17]), .IN3(core_block[49]), .IN4(n1128), .Q(
          n677));
   AO22X1 U697 (.IN1(n1060), .IN2(write_data[18]), .IN3(core_block[50]), .IN4(n1128), .Q(
          n678));
   AO22X1 U698 (.IN1(n1060), .IN2(write_data[19]), .IN3(core_block[51]), .IN4(n1128), .Q(
          n679));
   AO22X1 U699 (.IN1(n1060), .IN2(write_data[20]), .IN3(core_block[52]), .IN4(n1127), .Q(
          n680));
   AO22X1 U700 (.IN1(n1060), .IN2(write_data[21]), .IN3(core_block[53]), .IN4(n1127), .Q(
          n681));
   AO22X1 U701 (.IN1(n1060), .IN2(write_data[22]), .IN3(core_block[54]), .IN4(n1127), .Q(
          n682));
   AO22X1 U702 (.IN1(n1060), .IN2(write_data[23]), .IN3(core_block[55]), .IN4(n1127), .Q(
          n683));
   AO22X1 U703 (.IN1(n1061), .IN2(write_data[24]), .IN3(core_block[56]), .IN4(n1127), .Q(
          n684));
   AO22X1 U704 (.IN1(n1061), .IN2(write_data[25]), .IN3(core_block[57]), .IN4(n1127), .Q(
          n685));
   AO22X1 U705 (.IN1(n1061), .IN2(write_data[26]), .IN3(core_block[58]), .IN4(n1127), .Q(
          n686));
   AO22X1 U706 (.IN1(n1061), .IN2(write_data[27]), .IN3(core_block[59]), .IN4(n1127), .Q(
          n687));
   AO22X1 U707 (.IN1(n1061), .IN2(write_data[28]), .IN3(core_block[60]), .IN4(n1127), .Q(
          n688));
   AO22X1 U708 (.IN1(n1061), .IN2(write_data[29]), .IN3(core_block[61]), .IN4(n1127), .Q(
          n689));
   AO22X1 U709 (.IN1(n1061), .IN2(write_data[30]), .IN3(core_block[62]), .IN4(n1127), .Q(
          n690));
   AO22X1 U710 (.IN1(n1061), .IN2(write_data[31]), .IN3(core_block[63]), .IN4(n1127), .Q(
          n691));
   AO22X1 U711 (.IN1(n1056), .IN2(write_data[0]), .IN3(core_block[64]), .IN4(n612), .Q(
          n692));
   AO22X1 U712 (.IN1(n1056), .IN2(write_data[1]), .IN3(core_block[65]), .IN4(n612), .Q(
          n693));
   AO22X1 U713 (.IN1(n1056), .IN2(write_data[2]), .IN3(core_block[66]), .IN4(n612), .Q(
          n694));
   AO22X1 U714 (.IN1(n1056), .IN2(write_data[3]), .IN3(core_block[67]), .IN4(n612), .Q(
          n695));
   AO22X1 U715 (.IN1(n1056), .IN2(write_data[4]), .IN3(core_block[68]), .IN4(n612), .Q(
          n696));
   AO22X1 U716 (.IN1(n1056), .IN2(write_data[5]), .IN3(core_block[69]), .IN4(n612), .Q(
          n697));
   AO22X1 U717 (.IN1(n1056), .IN2(write_data[6]), .IN3(core_block[70]), .IN4(n612), .Q(
          n698));
   AO22X1 U718 (.IN1(n1056), .IN2(write_data[7]), .IN3(core_block[71]), .IN4(n612), .Q(
          n699));
   AO22X1 U719 (.IN1(n1056), .IN2(write_data[8]), .IN3(core_block[72]), .IN4(n1126), .Q(
          n700));
   AO22X1 U720 (.IN1(n1056), .IN2(write_data[9]), .IN3(core_block[73]), .IN4(n1126), .Q(
          n701));
   AO22X1 U721 (.IN1(n1056), .IN2(write_data[10]), .IN3(core_block[74]), .IN4(n1126), .Q(
          n702));
   AO22X1 U722 (.IN1(n1056), .IN2(write_data[11]), .IN3(core_block[75]), .IN4(n1126), .Q(
          n703));
   AO22X1 U723 (.IN1(n1057), .IN2(write_data[12]), .IN3(core_block[76]), .IN4(n1126), .Q(
          n704));
   AO22X1 U724 (.IN1(n1057), .IN2(write_data[13]), .IN3(core_block[77]), .IN4(n1126), .Q(
          n705));
   AO22X1 U725 (.IN1(n1057), .IN2(write_data[14]), .IN3(core_block[78]), .IN4(n1126), .Q(
          n706));
   AO22X1 U726 (.IN1(n1057), .IN2(write_data[15]), .IN3(core_block[79]), .IN4(n1126), .Q(
          n707));
   AO22X1 U727 (.IN1(n1057), .IN2(write_data[16]), .IN3(core_block[80]), .IN4(n1126), .Q(
          n708));
   AO22X1 U728 (.IN1(n1057), .IN2(write_data[17]), .IN3(core_block[81]), .IN4(n1126), .Q(
          n709));
   AO22X1 U729 (.IN1(n1057), .IN2(write_data[18]), .IN3(core_block[82]), .IN4(n1126), .Q(
          n710));
   AO22X1 U730 (.IN1(n1057), .IN2(write_data[19]), .IN3(core_block[83]), .IN4(n1126), .Q(
          n711));
   AO22X1 U731 (.IN1(n1057), .IN2(write_data[20]), .IN3(core_block[84]), .IN4(n1125), .Q(
          n712));
   AO22X1 U732 (.IN1(n1057), .IN2(write_data[21]), .IN3(core_block[85]), .IN4(n1125), .Q(
          n713));
   AO22X1 U733 (.IN1(n1057), .IN2(write_data[22]), .IN3(core_block[86]), .IN4(n1125), .Q(
          n714));
   AO22X1 U734 (.IN1(n1057), .IN2(write_data[23]), .IN3(core_block[87]), .IN4(n1125), .Q(
          n715));
   AO22X1 U735 (.IN1(n1058), .IN2(write_data[24]), .IN3(core_block[88]), .IN4(n1125), .Q(
          n716));
   AO22X1 U736 (.IN1(n1058), .IN2(write_data[25]), .IN3(core_block[89]), .IN4(n1125), .Q(
          n717));
   AO22X1 U737 (.IN1(n1058), .IN2(write_data[26]), .IN3(core_block[90]), .IN4(n1125), .Q(
          n718));
   AO22X1 U738 (.IN1(n1058), .IN2(write_data[27]), .IN3(core_block[91]), .IN4(n1125), .Q(
          n719));
   AO22X1 U739 (.IN1(n1058), .IN2(write_data[28]), .IN3(core_block[92]), .IN4(n1125), .Q(
          n720));
   AO22X1 U740 (.IN1(n1058), .IN2(write_data[29]), .IN3(core_block[93]), .IN4(n1125), .Q(
          n721));
   AO22X1 U741 (.IN1(n1058), .IN2(write_data[30]), .IN3(core_block[94]), .IN4(n1125), .Q(
          n722));
   AO22X1 U742 (.IN1(n1058), .IN2(write_data[31]), .IN3(core_block[95]), .IN4(n1125), .Q(
          n723));
   AO22X1 U743 (.IN1(n1053), .IN2(write_data[0]), .IN3(core_block[96]), .IN4(n613), .Q(
          n724));
   AO22X1 U744 (.IN1(n1053), .IN2(write_data[1]), .IN3(core_block[97]), .IN4(n613), .Q(
          n725));
   AO22X1 U745 (.IN1(n1053), .IN2(write_data[2]), .IN3(core_block[98]), .IN4(n613), .Q(
          n726));
   AO22X1 U746 (.IN1(n1053), .IN2(write_data[3]), .IN3(core_block[99]), .IN4(n613), .Q(
          n727));
   AO22X1 U747 (.IN1(n1053), .IN2(write_data[4]), .IN3(core_block[100]), .IN4(n613), .Q(
          n728));
   AO22X1 U748 (.IN1(n1053), .IN2(write_data[5]), .IN3(core_block[101]), .IN4(n613), .Q(
          n729));
   AO22X1 U749 (.IN1(n1053), .IN2(write_data[6]), .IN3(core_block[102]), .IN4(n613), .Q(
          n730));
   AO22X1 U750 (.IN1(n1053), .IN2(write_data[7]), .IN3(core_block[103]), .IN4(n613), .Q(
          n731));
   AO22X1 U751 (.IN1(n1053), .IN2(write_data[8]), .IN3(core_block[104]), .IN4(n1124), .Q(
          n732));
   AO22X1 U752 (.IN1(n1053), .IN2(write_data[9]), .IN3(core_block[105]), .IN4(n1124), .Q(
          n733));
   AO22X1 U753 (.IN1(n1053), .IN2(write_data[10]), .IN3(core_block[106]), .IN4(n1124), .Q(
          n734));
   AO22X1 U754 (.IN1(n1053), .IN2(write_data[11]), .IN3(core_block[107]), .IN4(n1124), .Q(
          n735));
   AO22X1 U755 (.IN1(n1054), .IN2(write_data[12]), .IN3(core_block[108]), .IN4(n1124), .Q(
          n736));
   AO22X1 U756 (.IN1(n1054), .IN2(write_data[13]), .IN3(core_block[109]), .IN4(n1124), .Q(
          n737));
   AO22X1 U757 (.IN1(n1054), .IN2(write_data[14]), .IN3(core_block[110]), .IN4(n1124), .Q(
          n738));
   AO22X1 U758 (.IN1(n1054), .IN2(write_data[15]), .IN3(core_block[111]), .IN4(n1124), .Q(
          n739));
   AO22X1 U759 (.IN1(n1054), .IN2(write_data[16]), .IN3(core_block[112]), .IN4(n1124), .Q(
          n740));
   AO22X1 U760 (.IN1(n1054), .IN2(write_data[17]), .IN3(core_block[113]), .IN4(n1124), .Q(
          n741));
   AO22X1 U761 (.IN1(n1054), .IN2(write_data[18]), .IN3(core_block[114]), .IN4(n1124), .Q(
          n742));
   AO22X1 U762 (.IN1(n1054), .IN2(write_data[19]), .IN3(core_block[115]), .IN4(n1124), .Q(
          n743));
   AO22X1 U763 (.IN1(n1054), .IN2(write_data[20]), .IN3(core_block[116]), .IN4(n1123), .Q(
          n744));
   AO22X1 U764 (.IN1(n1054), .IN2(write_data[21]), .IN3(core_block[117]), .IN4(n1123), .Q(
          n745));
   AO22X1 U765 (.IN1(n1054), .IN2(write_data[22]), .IN3(core_block[118]), .IN4(n1123), .Q(
          n746));
   AO22X1 U766 (.IN1(n1054), .IN2(write_data[23]), .IN3(core_block[119]), .IN4(n1123), .Q(
          n747));
   AO22X1 U767 (.IN1(n1055), .IN2(write_data[24]), .IN3(core_block[120]), .IN4(n1123), .Q(
          n748));
   AO22X1 U768 (.IN1(n1055), .IN2(write_data[25]), .IN3(core_block[121]), .IN4(n1123), .Q(
          n749));
   AO22X1 U769 (.IN1(n1055), .IN2(write_data[26]), .IN3(core_block[122]), .IN4(n1123), .Q(
          n750));
   AO22X1 U770 (.IN1(n1055), .IN2(write_data[27]), .IN3(core_block[123]), .IN4(n1123), .Q(
          n751));
   AO22X1 U771 (.IN1(n1055), .IN2(write_data[28]), .IN3(core_block[124]), .IN4(n1123), .Q(
          n752));
   AO22X1 U772 (.IN1(n1055), .IN2(write_data[29]), .IN3(core_block[125]), .IN4(n1123), .Q(
          n753));
   AO22X1 U773 (.IN1(n1055), .IN2(write_data[30]), .IN3(core_block[126]), .IN4(n1123), .Q(
          n754));
   AO22X1 U774 (.IN1(n1055), .IN2(write_data[31]), .IN3(core_block[127]), .IN4(n1123), .Q(
          n755));
   AND3X1 U775 (.IN1(n606), .IN2(n615), .IN3(N64), .Q(n608));
   NAND4X0 U778 (.IN1(n606), .IN2(address[3]), .IN3(n611), .IN4(n592), .QN(n616));
   AO22X1 U779 (.IN1(n1050), .IN2(write_data[0]), .IN3(core_key[0]), .IN4(n617), .Q(n758)
          );
   AO22X1 U780 (.IN1(n1050), .IN2(write_data[1]), .IN3(core_key[1]), .IN4(n617), .Q(n759)
          );
   AO22X1 U781 (.IN1(n1050), .IN2(write_data[2]), .IN3(core_key[2]), .IN4(n617), .Q(n760)
          );
   AO22X1 U782 (.IN1(n1050), .IN2(write_data[3]), .IN3(core_key[3]), .IN4(n617), .Q(n761)
          );
   AO22X1 U783 (.IN1(n1050), .IN2(write_data[4]), .IN3(core_key[4]), .IN4(n617), .Q(n762)
          );
   AO22X1 U784 (.IN1(n1050), .IN2(write_data[5]), .IN3(core_key[5]), .IN4(n617), .Q(n763)
          );
   AO22X1 U785 (.IN1(n1050), .IN2(write_data[6]), .IN3(core_key[6]), .IN4(n617), .Q(n764)
          );
   AO22X1 U786 (.IN1(n1050), .IN2(write_data[7]), .IN3(core_key[7]), .IN4(n617), .Q(n765)
          );
   AO22X1 U787 (.IN1(n1050), .IN2(write_data[8]), .IN3(core_key[8]), .IN4(n1122), .Q(n766)
          );
   AO22X1 U788 (.IN1(n1050), .IN2(write_data[9]), .IN3(core_key[9]), .IN4(n1122), .Q(n767)
          );
   AO22X1 U789 (.IN1(n1050), .IN2(write_data[10]), .IN3(core_key[10]), .IN4(n1122), .Q(
          n768));
   AO22X1 U790 (.IN1(n1050), .IN2(write_data[11]), .IN3(core_key[11]), .IN4(n1122), .Q(
          n769));
   AO22X1 U791 (.IN1(n1051), .IN2(write_data[12]), .IN3(core_key[12]), .IN4(n1122), .Q(
          n770));
   AO22X1 U792 (.IN1(n1051), .IN2(write_data[13]), .IN3(core_key[13]), .IN4(n1122), .Q(
          n771));
   AO22X1 U793 (.IN1(n1051), .IN2(write_data[14]), .IN3(core_key[14]), .IN4(n1122), .Q(
          n772));
   AO22X1 U794 (.IN1(n1051), .IN2(write_data[15]), .IN3(core_key[15]), .IN4(n1122), .Q(
          n773));
   AO22X1 U795 (.IN1(n1051), .IN2(write_data[16]), .IN3(core_key[16]), .IN4(n1122), .Q(
          n774));
   AO22X1 U796 (.IN1(n1051), .IN2(write_data[17]), .IN3(core_key[17]), .IN4(n1122), .Q(
          n775));
   AO22X1 U797 (.IN1(n1051), .IN2(write_data[18]), .IN3(core_key[18]), .IN4(n1122), .Q(
          n776));
   AO22X1 U798 (.IN1(n1051), .IN2(write_data[19]), .IN3(core_key[19]), .IN4(n1122), .Q(
          n777));
   AO22X1 U799 (.IN1(n1051), .IN2(write_data[20]), .IN3(core_key[20]), .IN4(n1121), .Q(
          n778));
   AO22X1 U800 (.IN1(n1051), .IN2(write_data[21]), .IN3(core_key[21]), .IN4(n1121), .Q(
          n779));
   AO22X1 U801 (.IN1(n1051), .IN2(write_data[22]), .IN3(core_key[22]), .IN4(n1121), .Q(
          n780));
   AO22X1 U802 (.IN1(n1051), .IN2(write_data[23]), .IN3(core_key[23]), .IN4(n1121), .Q(
          n781));
   AO22X1 U803 (.IN1(n1052), .IN2(write_data[24]), .IN3(core_key[24]), .IN4(n1121), .Q(
          n782));
   AO22X1 U804 (.IN1(n1052), .IN2(write_data[25]), .IN3(core_key[25]), .IN4(n1121), .Q(
          n783));
   AO22X1 U805 (.IN1(n1052), .IN2(write_data[26]), .IN3(core_key[26]), .IN4(n1121), .Q(
          n784));
   AO22X1 U806 (.IN1(n1052), .IN2(write_data[27]), .IN3(core_key[27]), .IN4(n1121), .Q(
          n785));
   AO22X1 U807 (.IN1(n1052), .IN2(write_data[28]), .IN3(core_key[28]), .IN4(n1121), .Q(
          n786));
   AO22X1 U808 (.IN1(n1052), .IN2(write_data[29]), .IN3(core_key[29]), .IN4(n1121), .Q(
          n787));
   AO22X1 U809 (.IN1(n1052), .IN2(write_data[30]), .IN3(core_key[30]), .IN4(n1121), .Q(
          n788));
   AO22X1 U810 (.IN1(n1052), .IN2(write_data[31]), .IN3(core_key[31]), .IN4(n1121), .Q(
          n789));
   AO22X1 U811 (.IN1(n1047), .IN2(write_data[0]), .IN3(core_key[32]), .IN4(n619), .Q(n790)
          );
   AO22X1 U812 (.IN1(n1047), .IN2(write_data[1]), .IN3(core_key[33]), .IN4(n619), .Q(n791)
          );
   AO22X1 U813 (.IN1(n1047), .IN2(write_data[2]), .IN3(core_key[34]), .IN4(n619), .Q(n792)
          );
   AO22X1 U814 (.IN1(n1047), .IN2(write_data[3]), .IN3(core_key[35]), .IN4(n619), .Q(n793)
          );
   AO22X1 U815 (.IN1(n1047), .IN2(write_data[4]), .IN3(core_key[36]), .IN4(n619), .Q(n794)
          );
   AO22X1 U816 (.IN1(n1047), .IN2(write_data[5]), .IN3(core_key[37]), .IN4(n619), .Q(n795)
          );
   AO22X1 U817 (.IN1(n1047), .IN2(write_data[6]), .IN3(core_key[38]), .IN4(n619), .Q(n796)
          );
   AO22X1 U818 (.IN1(n1047), .IN2(write_data[7]), .IN3(core_key[39]), .IN4(n619), .Q(n797)
          );
   AO22X1 U819 (.IN1(n1047), .IN2(write_data[8]), .IN3(core_key[40]), .IN4(n1120), .Q(n798)
          );
   AO22X1 U820 (.IN1(n1047), .IN2(write_data[9]), .IN3(core_key[41]), .IN4(n1120), .Q(n799)
          );
   AO22X1 U821 (.IN1(n1047), .IN2(write_data[10]), .IN3(core_key[42]), .IN4(n1120), .Q(
          n800));
   AO22X1 U822 (.IN1(n1047), .IN2(write_data[11]), .IN3(core_key[43]), .IN4(n1120), .Q(
          n801));
   AO22X1 U823 (.IN1(n1048), .IN2(write_data[12]), .IN3(core_key[44]), .IN4(n1120), .Q(
          n802));
   AO22X1 U824 (.IN1(n1048), .IN2(write_data[13]), .IN3(core_key[45]), .IN4(n1120), .Q(
          n803));
   AO22X1 U825 (.IN1(n1048), .IN2(write_data[14]), .IN3(core_key[46]), .IN4(n1120), .Q(
          n804));
   AO22X1 U826 (.IN1(n1048), .IN2(write_data[15]), .IN3(core_key[47]), .IN4(n1120), .Q(
          n805));
   AO22X1 U827 (.IN1(n1048), .IN2(write_data[16]), .IN3(core_key[48]), .IN4(n1120), .Q(
          n806));
   AO22X1 U828 (.IN1(n1048), .IN2(write_data[17]), .IN3(core_key[49]), .IN4(n1120), .Q(
          n807));
   AO22X1 U829 (.IN1(n1048), .IN2(write_data[18]), .IN3(core_key[50]), .IN4(n1120), .Q(
          n808));
   AO22X1 U830 (.IN1(n1048), .IN2(write_data[19]), .IN3(core_key[51]), .IN4(n1120), .Q(
          n809));
   AO22X1 U831 (.IN1(n1048), .IN2(write_data[20]), .IN3(core_key[52]), .IN4(n1119), .Q(
          n810));
   AO22X1 U832 (.IN1(n1048), .IN2(write_data[21]), .IN3(core_key[53]), .IN4(n1119), .Q(
          n811));
   AO22X1 U833 (.IN1(n1048), .IN2(write_data[22]), .IN3(core_key[54]), .IN4(n1119), .Q(
          n812));
   AO22X1 U834 (.IN1(n1048), .IN2(write_data[23]), .IN3(core_key[55]), .IN4(n1119), .Q(
          n813));
   AO22X1 U835 (.IN1(n1049), .IN2(write_data[24]), .IN3(core_key[56]), .IN4(n1119), .Q(
          n814));
   AO22X1 U836 (.IN1(n1049), .IN2(write_data[25]), .IN3(core_key[57]), .IN4(n1119), .Q(
          n815));
   AO22X1 U837 (.IN1(n1049), .IN2(write_data[26]), .IN3(core_key[58]), .IN4(n1119), .Q(
          n816));
   AO22X1 U838 (.IN1(n1049), .IN2(write_data[27]), .IN3(core_key[59]), .IN4(n1119), .Q(
          n817));
   AO22X1 U839 (.IN1(n1049), .IN2(write_data[28]), .IN3(core_key[60]), .IN4(n1119), .Q(
          n818));
   AO22X1 U840 (.IN1(n1049), .IN2(write_data[29]), .IN3(core_key[61]), .IN4(n1119), .Q(
          n819));
   AO22X1 U841 (.IN1(n1049), .IN2(write_data[30]), .IN3(core_key[62]), .IN4(n1119), .Q(
          n820));
   AO22X1 U842 (.IN1(n1049), .IN2(write_data[31]), .IN3(core_key[63]), .IN4(n1119), .Q(
          n821));
   AO22X1 U843 (.IN1(n1044), .IN2(write_data[0]), .IN3(core_key[64]), .IN4(n620), .Q(n822)
          );
   AO22X1 U844 (.IN1(n1044), .IN2(write_data[1]), .IN3(core_key[65]), .IN4(n620), .Q(n823)
          );
   AO22X1 U845 (.IN1(n1044), .IN2(write_data[2]), .IN3(core_key[66]), .IN4(n620), .Q(n824)
          );
   AO22X1 U846 (.IN1(n1044), .IN2(write_data[3]), .IN3(core_key[67]), .IN4(n620), .Q(n825)
          );
   AO22X1 U847 (.IN1(n1044), .IN2(write_data[4]), .IN3(core_key[68]), .IN4(n620), .Q(n826)
          );
   AO22X1 U848 (.IN1(n1044), .IN2(write_data[5]), .IN3(core_key[69]), .IN4(n620), .Q(n827)
          );
   AO22X1 U849 (.IN1(n1044), .IN2(write_data[6]), .IN3(core_key[70]), .IN4(n620), .Q(n828)
          );
   AO22X1 U850 (.IN1(n1044), .IN2(write_data[7]), .IN3(core_key[71]), .IN4(n620), .Q(n829)
          );
   AO22X1 U851 (.IN1(n1044), .IN2(write_data[8]), .IN3(core_key[72]), .IN4(n1118), .Q(n830)
          );
   AO22X1 U852 (.IN1(n1044), .IN2(write_data[9]), .IN3(core_key[73]), .IN4(n1118), .Q(n831)
          );
   AO22X1 U853 (.IN1(n1044), .IN2(write_data[10]), .IN3(core_key[74]), .IN4(n1118), .Q(
          n832));
   AO22X1 U854 (.IN1(n1044), .IN2(write_data[11]), .IN3(core_key[75]), .IN4(n1118), .Q(
          n833));
   AO22X1 U855 (.IN1(n1045), .IN2(write_data[12]), .IN3(core_key[76]), .IN4(n1118), .Q(
          n834));
   AO22X1 U856 (.IN1(n1045), .IN2(write_data[13]), .IN3(core_key[77]), .IN4(n1118), .Q(
          n835));
   AO22X1 U857 (.IN1(n1045), .IN2(write_data[14]), .IN3(core_key[78]), .IN4(n1118), .Q(
          n836));
   AO22X1 U858 (.IN1(n1045), .IN2(write_data[15]), .IN3(core_key[79]), .IN4(n1118), .Q(
          n837));
   AO22X1 U859 (.IN1(n1045), .IN2(write_data[16]), .IN3(core_key[80]), .IN4(n1118), .Q(
          n838));
   AO22X1 U860 (.IN1(n1045), .IN2(write_data[17]), .IN3(core_key[81]), .IN4(n1118), .Q(
          n839));
   AO22X1 U861 (.IN1(n1045), .IN2(write_data[18]), .IN3(core_key[82]), .IN4(n1118), .Q(
          n840));
   AO22X1 U862 (.IN1(n1045), .IN2(write_data[19]), .IN3(core_key[83]), .IN4(n1118), .Q(
          n841));
   AO22X1 U863 (.IN1(n1045), .IN2(write_data[20]), .IN3(core_key[84]), .IN4(n1117), .Q(
          n842));
   AO22X1 U864 (.IN1(n1045), .IN2(write_data[21]), .IN3(core_key[85]), .IN4(n1117), .Q(
          n843));
   AO22X1 U865 (.IN1(n1045), .IN2(write_data[22]), .IN3(core_key[86]), .IN4(n1117), .Q(
          n844));
   AO22X1 U866 (.IN1(n1045), .IN2(write_data[23]), .IN3(core_key[87]), .IN4(n1117), .Q(
          n845));
   AO22X1 U867 (.IN1(n1046), .IN2(write_data[24]), .IN3(core_key[88]), .IN4(n1117), .Q(
          n846));
   AO22X1 U868 (.IN1(n1046), .IN2(write_data[25]), .IN3(core_key[89]), .IN4(n1117), .Q(
          n847));
   AO22X1 U869 (.IN1(n1046), .IN2(write_data[26]), .IN3(core_key[90]), .IN4(n1117), .Q(
          n848));
   AO22X1 U870 (.IN1(n1046), .IN2(write_data[27]), .IN3(core_key[91]), .IN4(n1117), .Q(
          n849));
   AO22X1 U871 (.IN1(n1046), .IN2(write_data[28]), .IN3(core_key[92]), .IN4(n1117), .Q(
          n850));
   AO22X1 U872 (.IN1(n1046), .IN2(write_data[29]), .IN3(core_key[93]), .IN4(n1117), .Q(
          n851));
   AO22X1 U873 (.IN1(n1046), .IN2(write_data[30]), .IN3(core_key[94]), .IN4(n1117), .Q(
          n852));
   AO22X1 U874 (.IN1(n1046), .IN2(write_data[31]), .IN3(core_key[95]), .IN4(n1117), .Q(
          n853));
   AO22X1 U875 (.IN1(n1041), .IN2(write_data[0]), .IN3(core_key[96]), .IN4(n621), .Q(n854)
          );
   AO22X1 U876 (.IN1(n1041), .IN2(write_data[1]), .IN3(core_key[97]), .IN4(n621), .Q(n855)
          );
   AO22X1 U877 (.IN1(n1041), .IN2(write_data[2]), .IN3(core_key[98]), .IN4(n621), .Q(n856)
          );
   AO22X1 U878 (.IN1(n1041), .IN2(write_data[3]), .IN3(core_key[99]), .IN4(n621), .Q(n857)
          );
   AO22X1 U879 (.IN1(n1041), .IN2(write_data[4]), .IN3(core_key[100]), .IN4(n621), .Q(n858)
          );
   AO22X1 U880 (.IN1(n1041), .IN2(write_data[5]), .IN3(core_key[101]), .IN4(n621), .Q(n859)
          );
   AO22X1 U881 (.IN1(n1041), .IN2(write_data[6]), .IN3(core_key[102]), .IN4(n621), .Q(n860)
          );
   AO22X1 U882 (.IN1(n1041), .IN2(write_data[7]), .IN3(core_key[103]), .IN4(n621), .Q(n861)
          );
   AO22X1 U883 (.IN1(n1041), .IN2(write_data[8]), .IN3(core_key[104]), .IN4(n1116), .Q(
          n862));
   AO22X1 U884 (.IN1(n1041), .IN2(write_data[9]), .IN3(core_key[105]), .IN4(n1116), .Q(
          n863));
   AO22X1 U885 (.IN1(n1041), .IN2(write_data[10]), .IN3(core_key[106]), .IN4(n1116), .Q(
          n864));
   AO22X1 U886 (.IN1(n1041), .IN2(write_data[11]), .IN3(core_key[107]), .IN4(n1116), .Q(
          n865));
   AO22X1 U887 (.IN1(n1042), .IN2(write_data[12]), .IN3(core_key[108]), .IN4(n1116), .Q(
          n866));
   AO22X1 U888 (.IN1(n1042), .IN2(write_data[13]), .IN3(core_key[109]), .IN4(n1116), .Q(
          n867));
   AO22X1 U889 (.IN1(n1042), .IN2(write_data[14]), .IN3(core_key[110]), .IN4(n1116), .Q(
          n868));
   AO22X1 U890 (.IN1(n1042), .IN2(write_data[15]), .IN3(core_key[111]), .IN4(n1116), .Q(
          n869));
   AO22X1 U891 (.IN1(n1042), .IN2(write_data[16]), .IN3(core_key[112]), .IN4(n1116), .Q(
          n870));
   AO22X1 U892 (.IN1(n1042), .IN2(write_data[17]), .IN3(core_key[113]), .IN4(n1116), .Q(
          n871));
   AO22X1 U893 (.IN1(n1042), .IN2(write_data[18]), .IN3(core_key[114]), .IN4(n1116), .Q(
          n872));
   AO22X1 U894 (.IN1(n1042), .IN2(write_data[19]), .IN3(core_key[115]), .IN4(n1116), .Q(
          n873));
   AO22X1 U895 (.IN1(n1042), .IN2(write_data[20]), .IN3(core_key[116]), .IN4(n1115), .Q(
          n874));
   AO22X1 U896 (.IN1(n1042), .IN2(write_data[21]), .IN3(core_key[117]), .IN4(n1115), .Q(
          n875));
   AO22X1 U897 (.IN1(n1042), .IN2(write_data[22]), .IN3(core_key[118]), .IN4(n1115), .Q(
          n876));
   AO22X1 U898 (.IN1(n1042), .IN2(write_data[23]), .IN3(core_key[119]), .IN4(n1115), .Q(
          n877));
   AO22X1 U899 (.IN1(n1043), .IN2(write_data[24]), .IN3(core_key[120]), .IN4(n1115), .Q(
          n878));
   AO22X1 U900 (.IN1(n1043), .IN2(write_data[25]), .IN3(core_key[121]), .IN4(n1115), .Q(
          n879));
   AO22X1 U901 (.IN1(n1043), .IN2(write_data[26]), .IN3(core_key[122]), .IN4(n1115), .Q(
          n880));
   AO22X1 U902 (.IN1(n1043), .IN2(write_data[27]), .IN3(core_key[123]), .IN4(n1115), .Q(
          n881));
   AO22X1 U903 (.IN1(n1043), .IN2(write_data[28]), .IN3(core_key[124]), .IN4(n1115), .Q(
          n882));
   AO22X1 U904 (.IN1(n1043), .IN2(write_data[29]), .IN3(core_key[125]), .IN4(n1115), .Q(
          n883));
   AO22X1 U905 (.IN1(n1043), .IN2(write_data[30]), .IN3(core_key[126]), .IN4(n1115), .Q(
          n884));
   AO22X1 U906 (.IN1(n1043), .IN2(write_data[31]), .IN3(core_key[127]), .IN4(n1115), .Q(
          n885));
   AND2X1 U907 (.IN1(address[2]), .IN2(n622), .Q(n618));
   AO22X1 U908 (.IN1(n1038), .IN2(write_data[0]), .IN3(core_key[128]), .IN4(n623), .Q(n886)
          );
   AO22X1 U909 (.IN1(n1038), .IN2(write_data[1]), .IN3(core_key[129]), .IN4(n623), .Q(n887)
          );
   AO22X1 U910 (.IN1(n1038), .IN2(write_data[2]), .IN3(core_key[130]), .IN4(n623), .Q(n888)
          );
   AO22X1 U911 (.IN1(n1038), .IN2(write_data[3]), .IN3(core_key[131]), .IN4(n623), .Q(n889)
          );
   AO22X1 U912 (.IN1(n1038), .IN2(write_data[4]), .IN3(core_key[132]), .IN4(n623), .Q(n890)
          );
   AO22X1 U913 (.IN1(n1038), .IN2(write_data[5]), .IN3(core_key[133]), .IN4(n623), .Q(n891)
          );
   AO22X1 U914 (.IN1(n1038), .IN2(write_data[6]), .IN3(core_key[134]), .IN4(n623), .Q(n892)
          );
   AO22X1 U915 (.IN1(n1038), .IN2(write_data[7]), .IN3(core_key[135]), .IN4(n623), .Q(n893)
          );
   AO22X1 U916 (.IN1(n1038), .IN2(write_data[8]), .IN3(core_key[136]), .IN4(n1114), .Q(
          n894));
   AO22X1 U917 (.IN1(n1038), .IN2(write_data[9]), .IN3(core_key[137]), .IN4(n1114), .Q(
          n895));
   AO22X1 U918 (.IN1(n1038), .IN2(write_data[10]), .IN3(core_key[138]), .IN4(n1114), .Q(
          n896));
   AO22X1 U919 (.IN1(n1038), .IN2(write_data[11]), .IN3(core_key[139]), .IN4(n1114), .Q(
          n897));
   AO22X1 U920 (.IN1(n1039), .IN2(write_data[12]), .IN3(core_key[140]), .IN4(n1114), .Q(
          n898));
   AO22X1 U921 (.IN1(n1039), .IN2(write_data[13]), .IN3(core_key[141]), .IN4(n1114), .Q(
          n899));
   AO22X1 U922 (.IN1(n1039), .IN2(write_data[14]), .IN3(core_key[142]), .IN4(n1114), .Q(
          n900));
   AO22X1 U923 (.IN1(n1039), .IN2(write_data[15]), .IN3(core_key[143]), .IN4(n1114), .Q(
          n901));
   AO22X1 U924 (.IN1(n1039), .IN2(write_data[16]), .IN3(core_key[144]), .IN4(n1114), .Q(
          n902));
   AO22X1 U925 (.IN1(n1039), .IN2(write_data[17]), .IN3(core_key[145]), .IN4(n1114), .Q(
          n903));
   AO22X1 U926 (.IN1(n1039), .IN2(write_data[18]), .IN3(core_key[146]), .IN4(n1114), .Q(
          n904));
   AO22X1 U927 (.IN1(n1039), .IN2(write_data[19]), .IN3(core_key[147]), .IN4(n1114), .Q(
          n905));
   AO22X1 U928 (.IN1(n1039), .IN2(write_data[20]), .IN3(core_key[148]), .IN4(n1113), .Q(
          n906));
   AO22X1 U929 (.IN1(n1039), .IN2(write_data[21]), .IN3(core_key[149]), .IN4(n1113), .Q(
          n907));
   AO22X1 U930 (.IN1(n1039), .IN2(write_data[22]), .IN3(core_key[150]), .IN4(n1113), .Q(
          n908));
   AO22X1 U931 (.IN1(n1039), .IN2(write_data[23]), .IN3(core_key[151]), .IN4(n1113), .Q(
          n909));
   AO22X1 U932 (.IN1(n1040), .IN2(write_data[24]), .IN3(core_key[152]), .IN4(n1113), .Q(
          n910));
   AO22X1 U933 (.IN1(n1040), .IN2(write_data[25]), .IN3(core_key[153]), .IN4(n1113), .Q(
          n911));
   AO22X1 U934 (.IN1(n1040), .IN2(write_data[26]), .IN3(core_key[154]), .IN4(n1113), .Q(
          n912));
   AO22X1 U935 (.IN1(n1040), .IN2(write_data[27]), .IN3(core_key[155]), .IN4(n1113), .Q(
          n913));
   AO22X1 U936 (.IN1(n1040), .IN2(write_data[28]), .IN3(core_key[156]), .IN4(n1113), .Q(
          n914));
   AO22X1 U937 (.IN1(n1040), .IN2(write_data[29]), .IN3(core_key[157]), .IN4(n1113), .Q(
          n915));
   AO22X1 U938 (.IN1(n1040), .IN2(write_data[30]), .IN3(core_key[158]), .IN4(n1113), .Q(
          n916));
   AO22X1 U939 (.IN1(n1040), .IN2(write_data[31]), .IN3(core_key[159]), .IN4(n1113), .Q(
          n917));
   AND2X1 U940 (.IN1(n609), .IN2(n1159), .Q(n601));
   AO22X1 U941 (.IN1(n1035), .IN2(write_data[0]), .IN3(core_key[160]), .IN4(n624), .Q(n918)
          );
   AO22X1 U942 (.IN1(n1035), .IN2(write_data[1]), .IN3(core_key[161]), .IN4(n624), .Q(n919)
          );
   AO22X1 U943 (.IN1(n1035), .IN2(write_data[2]), .IN3(core_key[162]), .IN4(n624), .Q(n920)
          );
   AO22X1 U944 (.IN1(n1035), .IN2(write_data[3]), .IN3(core_key[163]), .IN4(n624), .Q(n921)
          );
   AO22X1 U945 (.IN1(n1035), .IN2(write_data[4]), .IN3(core_key[164]), .IN4(n624), .Q(n922)
          );
   AO22X1 U946 (.IN1(n1035), .IN2(write_data[5]), .IN3(core_key[165]), .IN4(n624), .Q(n923)
          );
   AO22X1 U947 (.IN1(n1035), .IN2(write_data[6]), .IN3(core_key[166]), .IN4(n624), .Q(n924)
          );
   AO22X1 U948 (.IN1(n1035), .IN2(write_data[7]), .IN3(core_key[167]), .IN4(n624), .Q(n925)
          );
   AO22X1 U949 (.IN1(n1035), .IN2(write_data[8]), .IN3(core_key[168]), .IN4(n1112), .Q(
          n926));
   AO22X1 U950 (.IN1(n1035), .IN2(write_data[9]), .IN3(core_key[169]), .IN4(n1112), .Q(
          n927));
   AO22X1 U951 (.IN1(n1035), .IN2(write_data[10]), .IN3(core_key[170]), .IN4(n1112), .Q(
          n928));
   AO22X1 U952 (.IN1(n1035), .IN2(write_data[11]), .IN3(core_key[171]), .IN4(n1112), .Q(
          n929));
   AO22X1 U953 (.IN1(n1036), .IN2(write_data[12]), .IN3(core_key[172]), .IN4(n1112), .Q(
          n930));
   AO22X1 U954 (.IN1(n1036), .IN2(write_data[13]), .IN3(core_key[173]), .IN4(n1112), .Q(
          n931));
   AO22X1 U955 (.IN1(n1036), .IN2(write_data[14]), .IN3(core_key[174]), .IN4(n1112), .Q(
          n932));
   AO22X1 U956 (.IN1(n1036), .IN2(write_data[15]), .IN3(core_key[175]), .IN4(n1112), .Q(
          n933));
   AO22X1 U957 (.IN1(n1036), .IN2(write_data[16]), .IN3(core_key[176]), .IN4(n1112), .Q(
          n934));
   AO22X1 U958 (.IN1(n1036), .IN2(write_data[17]), .IN3(core_key[177]), .IN4(n1112), .Q(
          n935));
   AO22X1 U959 (.IN1(n1036), .IN2(write_data[18]), .IN3(core_key[178]), .IN4(n1112), .Q(
          n936));
   AO22X1 U960 (.IN1(n1036), .IN2(write_data[19]), .IN3(core_key[179]), .IN4(n1112), .Q(
          n937));
   AO22X1 U961 (.IN1(n1036), .IN2(write_data[20]), .IN3(core_key[180]), .IN4(n1111), .Q(
          n938));
   AO22X1 U962 (.IN1(n1036), .IN2(write_data[21]), .IN3(core_key[181]), .IN4(n1111), .Q(
          n939));
   AO22X1 U963 (.IN1(n1036), .IN2(write_data[22]), .IN3(core_key[182]), .IN4(n1111), .Q(
          n940));
   AO22X1 U964 (.IN1(n1036), .IN2(write_data[23]), .IN3(core_key[183]), .IN4(n1111), .Q(
          n941));
   AO22X1 U965 (.IN1(n1037), .IN2(write_data[24]), .IN3(core_key[184]), .IN4(n1111), .Q(
          n942));
   AO22X1 U966 (.IN1(n1037), .IN2(write_data[25]), .IN3(core_key[185]), .IN4(n1111), .Q(
          n943));
   AO22X1 U967 (.IN1(n1037), .IN2(write_data[26]), .IN3(core_key[186]), .IN4(n1111), .Q(
          n944));
   AO22X1 U968 (.IN1(n1037), .IN2(write_data[27]), .IN3(core_key[187]), .IN4(n1111), .Q(
          n945));
   AO22X1 U969 (.IN1(n1037), .IN2(write_data[28]), .IN3(core_key[188]), .IN4(n1111), .Q(
          n946));
   AO22X1 U970 (.IN1(n1037), .IN2(write_data[29]), .IN3(core_key[189]), .IN4(n1111), .Q(
          n947));
   AO22X1 U971 (.IN1(n1037), .IN2(write_data[30]), .IN3(core_key[190]), .IN4(n1111), .Q(
          n948));
   AO22X1 U972 (.IN1(n1037), .IN2(write_data[31]), .IN3(core_key[191]), .IN4(n1111), .Q(
          n949));
   AND2X1 U973 (.IN1(n611), .IN2(n1159), .Q(n604));
   AO22X1 U974 (.IN1(n1032), .IN2(write_data[0]), .IN3(core_key[192]), .IN4(n625), .Q(n950)
          );
   AO22X1 U975 (.IN1(n1032), .IN2(write_data[1]), .IN3(core_key[193]), .IN4(n625), .Q(n951)
          );
   AO22X1 U976 (.IN1(n1032), .IN2(write_data[2]), .IN3(core_key[194]), .IN4(n625), .Q(n952)
          );
   AO22X1 U977 (.IN1(n1032), .IN2(write_data[3]), .IN3(core_key[195]), .IN4(n625), .Q(n953)
          );
   AO22X1 U978 (.IN1(n1032), .IN2(write_data[4]), .IN3(core_key[196]), .IN4(n625), .Q(n954)
          );
   AO22X1 U979 (.IN1(n1032), .IN2(write_data[5]), .IN3(core_key[197]), .IN4(n625), .Q(n955)
          );
   AO22X1 U980 (.IN1(n1032), .IN2(write_data[6]), .IN3(core_key[198]), .IN4(n625), .Q(n956)
          );
   AO22X1 U981 (.IN1(n1032), .IN2(write_data[7]), .IN3(core_key[199]), .IN4(n625), .Q(n957)
          );
   AO22X1 U982 (.IN1(n1032), .IN2(write_data[8]), .IN3(core_key[200]), .IN4(n1110), .Q(
          n958));
   AO22X1 U983 (.IN1(n1032), .IN2(write_data[9]), .IN3(core_key[201]), .IN4(n1110), .Q(
          n959));
   AO22X1 U984 (.IN1(n1032), .IN2(write_data[10]), .IN3(core_key[202]), .IN4(n1110), .Q(
          n960));
   AO22X1 U985 (.IN1(n1032), .IN2(write_data[11]), .IN3(core_key[203]), .IN4(n1110), .Q(
          n961));
   AO22X1 U986 (.IN1(n1033), .IN2(write_data[12]), .IN3(core_key[204]), .IN4(n1110), .Q(
          n962));
   AO22X1 U987 (.IN1(n1033), .IN2(write_data[13]), .IN3(core_key[205]), .IN4(n1110), .Q(
          n963));
   AO22X1 U988 (.IN1(n1033), .IN2(write_data[14]), .IN3(core_key[206]), .IN4(n1110), .Q(
          n964));
   AO22X1 U989 (.IN1(n1033), .IN2(write_data[15]), .IN3(core_key[207]), .IN4(n1110), .Q(
          n965));
   AO22X1 U990 (.IN1(n1033), .IN2(write_data[16]), .IN3(core_key[208]), .IN4(n1110), .Q(
          n966));
   AO22X1 U991 (.IN1(n1033), .IN2(write_data[17]), .IN3(core_key[209]), .IN4(n1110), .Q(
          n967));
   AO22X1 U992 (.IN1(n1033), .IN2(write_data[18]), .IN3(core_key[210]), .IN4(n1110), .Q(
          n968));
   AO22X1 U993 (.IN1(n1033), .IN2(write_data[19]), .IN3(core_key[211]), .IN4(n1110), .Q(
          n969));
   AO22X1 U994 (.IN1(n1033), .IN2(write_data[20]), .IN3(core_key[212]), .IN4(n1109), .Q(
          n970));
   AO22X1 U995 (.IN1(n1033), .IN2(write_data[21]), .IN3(core_key[213]), .IN4(n1109), .Q(
          n971));
   AO22X1 U996 (.IN1(n1033), .IN2(write_data[22]), .IN3(core_key[214]), .IN4(n1109), .Q(
          n972));
   AO22X1 U997 (.IN1(n1033), .IN2(write_data[23]), .IN3(core_key[215]), .IN4(n1109), .Q(
          n973));
   AO22X1 U998 (.IN1(n1034), .IN2(write_data[24]), .IN3(core_key[216]), .IN4(n1109), .Q(
          n974));
   AO22X1 U999 (.IN1(n1034), .IN2(write_data[25]), .IN3(core_key[217]), .IN4(n1109), .Q(
          n975));
   AO22X1 U1000 (.IN1(n1034), .IN2(write_data[26]), .IN3(core_key[218]), .IN4(n1109), .Q(
          n976));
   AO22X1 U1001 (.IN1(n1034), .IN2(write_data[27]), .IN3(core_key[219]), .IN4(n1109), .Q(
          n977));
   AO22X1 U1002 (.IN1(n1034), .IN2(write_data[28]), .IN3(core_key[220]), .IN4(n1109), .Q(
          n978));
   AO22X1 U1003 (.IN1(n1034), .IN2(write_data[29]), .IN3(core_key[221]), .IN4(n1109), .Q(
          n979));
   AO22X1 U1004 (.IN1(n1034), .IN2(write_data[30]), .IN3(core_key[222]), .IN4(n1109), .Q(
          n980));
   AO22X1 U1005 (.IN1(n1034), .IN2(write_data[31]), .IN3(core_key[223]), .IN4(n1109), .Q(
          n981));
   AND2X1 U1006 (.IN1(n598), .IN2(n1159), .Q(n603));
   AO22X1 U1007 (.IN1(n1029), .IN2(write_data[0]), .IN3(core_key[224]), .IN4(n626), .Q(
          n982));
   AO22X1 U1008 (.IN1(n1029), .IN2(write_data[1]), .IN3(core_key[225]), .IN4(n626), .Q(
          n983));
   AO22X1 U1009 (.IN1(n1029), .IN2(write_data[2]), .IN3(core_key[226]), .IN4(n626), .Q(
          n984));
   AO22X1 U1010 (.IN1(n1029), .IN2(write_data[3]), .IN3(core_key[227]), .IN4(n626), .Q(
          n985));
   AO22X1 U1011 (.IN1(n1029), .IN2(write_data[4]), .IN3(core_key[228]), .IN4(n626), .Q(
          n986));
   AO22X1 U1012 (.IN1(n1029), .IN2(write_data[5]), .IN3(core_key[229]), .IN4(n626), .Q(
          n987));
   AO22X1 U1013 (.IN1(n1029), .IN2(write_data[6]), .IN3(core_key[230]), .IN4(n626), .Q(
          n988));
   AO22X1 U1014 (.IN1(n1029), .IN2(write_data[7]), .IN3(core_key[231]), .IN4(n626), .Q(
          n989));
   AO22X1 U1015 (.IN1(n1029), .IN2(write_data[8]), .IN3(core_key[232]), .IN4(n1108), .Q(
          n990));
   AO22X1 U1016 (.IN1(n1029), .IN2(write_data[9]), .IN3(core_key[233]), .IN4(n1108), .Q(
          n991));
   AO22X1 U1017 (.IN1(n1029), .IN2(write_data[10]), .IN3(core_key[234]), .IN4(n1108), .Q(
          n992));
   AO22X1 U1018 (.IN1(n1029), .IN2(write_data[11]), .IN3(core_key[235]), .IN4(n1108), .Q(
          n993));
   AO22X1 U1019 (.IN1(n1030), .IN2(write_data[12]), .IN3(core_key[236]), .IN4(n1108), .Q(
          n994));
   AO22X1 U1020 (.IN1(n1030), .IN2(write_data[13]), .IN3(core_key[237]), .IN4(n1108), .Q(
          n995));
   AO22X1 U1021 (.IN1(n1030), .IN2(write_data[14]), .IN3(core_key[238]), .IN4(n1108), .Q(
          n996));
   AO22X1 U1022 (.IN1(n1030), .IN2(write_data[15]), .IN3(core_key[239]), .IN4(n1108), .Q(
          n997));
   AO22X1 U1023 (.IN1(n1030), .IN2(write_data[16]), .IN3(core_key[240]), .IN4(n1108), .Q(
          n998));
   AO22X1 U1024 (.IN1(n1030), .IN2(write_data[17]), .IN3(core_key[241]), .IN4(n1108), .Q(
          n999));
   AO22X1 U1025 (.IN1(n1030), .IN2(write_data[18]), .IN3(core_key[242]), .IN4(n1108), .Q(
          n1000));
   AO22X1 U1026 (.IN1(n1030), .IN2(write_data[19]), .IN3(core_key[243]), .IN4(n1108), .Q(
          n1001));
   AO22X1 U1027 (.IN1(n1030), .IN2(write_data[20]), .IN3(core_key[244]), .IN4(n1107), .Q(
          n1002));
   AO22X1 U1028 (.IN1(n1030), .IN2(write_data[21]), .IN3(core_key[245]), .IN4(n1107), .Q(
          n1003));
   AO22X1 U1029 (.IN1(n1030), .IN2(write_data[22]), .IN3(core_key[246]), .IN4(n1107), .Q(
          n1004));
   AO22X1 U1030 (.IN1(n1030), .IN2(write_data[23]), .IN3(core_key[247]), .IN4(n1107), .Q(
          n1005));
   AO22X1 U1031 (.IN1(n1031), .IN2(write_data[24]), .IN3(core_key[248]), .IN4(n1107), .Q(
          n1006));
   AO22X1 U1032 (.IN1(n1031), .IN2(write_data[25]), .IN3(core_key[249]), .IN4(n1107), .Q(
          n1007));
   AO22X1 U1033 (.IN1(n1031), .IN2(write_data[26]), .IN3(core_key[250]), .IN4(n1107), .Q(
          n1008));
   AO22X1 U1034 (.IN1(n1031), .IN2(write_data[27]), .IN3(core_key[251]), .IN4(n1107), .Q(
          n1009));
   AO22X1 U1035 (.IN1(n1031), .IN2(write_data[28]), .IN3(core_key[252]), .IN4(n1107), .Q(
          n1010));
   AO22X1 U1036 (.IN1(n1031), .IN2(write_data[29]), .IN3(core_key[253]), .IN4(n1107), .Q(
          n1011));
   AO22X1 U1037 (.IN1(n1031), .IN2(write_data[30]), .IN3(core_key[254]), .IN4(n1107), .Q(
          n1012));
   AO22X1 U1038 (.IN1(n1031), .IN2(write_data[31]), .IN3(core_key[255]), .IN4(n1107), .Q(
          n1013));
   AND2X1 U1039 (.IN1(n614), .IN2(n1159), .Q(n605));
   AND3X1 U1040 (.IN1(n606), .IN2(n627), .IN3(N62), .Q(n622));
   AND3X1 U1041 (.IN1(write_data[0]), .IN2(n1157), .IN3(n606), .Q(init_new));
   NAND3X0 U1042 (.IN1(n614), .IN2(n592), .IN3(address[3]), .QN(n599));
   OR2X1 U1043 (.IN1(address[4]), .IN2(n615), .Q(n627));
   OR3X1 U1044 (.IN1(address[7]), .IN2(address[6]), .IN3(address[5]), .Q(n615));
   aes_core_test_1 core (.clk(n1562_buf_net1), .reset_n(n1089), .encdec(core_encdec), .
          init(core_init), .next(core_next), .ready(core_ready), .key(core_key), .keylen(
          core_keylen), .block(core_block), .result(core_result), .result_valid(core_valid)
          , .test_si3(test_si4), .test_si2(TEST_SI3), .test_si1(n1429), .test_so3(n1422), .
          test_so2(TEST_SO3), .test_so1(TEST_SO1), .test_se(TEST_SE_buf_net1));
   NAND2X1 U1045 (.IN1(n618), .IN2(n614), .QN(n621));
   NAND2X1 U1046 (.IN1(n608), .IN2(n614), .QN(n613));
   NAND2X1 U1047 (.IN1(n618), .IN2(n611), .QN(n619));
   NAND2X1 U1048 (.IN1(n608), .IN2(n611), .QN(n610));
   NAND2X1 U1049 (.IN1(n618), .IN2(n598), .QN(n620));
   NAND2X1 U1050 (.IN1(n608), .IN2(n598), .QN(n612));
   NAND2X1 U1051 (.IN1(n618), .IN2(n609), .QN(n617));
   NAND2X1 U1052 (.IN1(n608), .IN2(n609), .QN(n607));
   NAND2X1 U1053 (.IN1(n604), .IN2(n602), .QN(n1014));
   NAND2X1 U1054 (.IN1(n601), .IN2(n602), .QN(n1015));
   NAND2X1 U1055 (.IN1(n605), .IN2(n602), .QN(n1016));
   NAND2X1 U1056 (.IN1(n603), .IN2(n602), .QN(n1017));
   NAND2X1 U1057 (.IN1(n622), .IN2(n605), .QN(n626));
   NAND2X1 U1058 (.IN1(n622), .IN2(n603), .QN(n625));
   NAND2X1 U1059 (.IN1(n622), .IN2(n604), .QN(n624));
   NAND2X1 U1060 (.IN1(n622), .IN2(n601), .QN(n623));
   NBUFFX2 U1061 (.INP(reset_n), .Z(n1143));
   NBUFFX2 U1062 (.INP(reset_n), .Z(n1144));
   NBUFFX2 U1063 (.INP(reset_n), .Z(n1145));
   NBUFFX2 U1064 (.INP(reset_n), .Z(n1146));
   NBUFFX2 U1065 (.INP(n1026), .Z(n1024));
   NBUFFX2 U1066 (.INP(n1026), .Z(n1023));
   NBUFFX2 U1067 (.INP(n1027), .Z(n1022));
   NBUFFX2 U1068 (.INP(n1027), .Z(n1021));
   NBUFFX2 U1069 (.INP(n1027), .Z(n1020));
   NBUFFX2 U1070 (.INP(n1028), .Z(n1019));
   NBUFFX2 U1071 (.INP(n1028), .Z(n1018));
   NBUFFX2 U1072 (.INP(n1026), .Z(n1025));
   INVX0 U1073 (.INP(n1064), .ZN(n1130));
   INVX0 U1074 (.INP(n1064), .ZN(n1129));
   INVX0 U1075 (.INP(n1061), .ZN(n1128));
   INVX0 U1076 (.INP(n1061), .ZN(n1127));
   INVX0 U1077 (.INP(n1055), .ZN(n1124));
   INVX0 U1078 (.INP(n1055), .ZN(n1123));
   INVX0 U1079 (.INP(n1052), .ZN(n1122));
   INVX0 U1080 (.INP(n1052), .ZN(n1121));
   INVX0 U1081 (.INP(n1049), .ZN(n1120));
   INVX0 U1082 (.INP(n1049), .ZN(n1119));
   INVX0 U1083 (.INP(n1043), .ZN(n1116));
   INVX0 U1084 (.INP(n1043), .ZN(n1115));
   INVX0 U1085 (.INP(n1058), .ZN(n1126));
   INVX0 U1086 (.INP(n1058), .ZN(n1125));
   INVX0 U1087 (.INP(n1046), .ZN(n1118));
   INVX0 U1088 (.INP(n1046), .ZN(n1117));
   INVX0 U1089 (.INP(n1040), .ZN(n1114));
   INVX0 U1090 (.INP(n1040), .ZN(n1113));
   INVX0 U1091 (.INP(n1037), .ZN(n1112));
   INVX0 U1092 (.INP(n1037), .ZN(n1111));
   INVX0 U1093 (.INP(n1034), .ZN(n1110));
   INVX0 U1094 (.INP(n1034), .ZN(n1109));
   INVX0 U1095 (.INP(n1031), .ZN(n1108));
   INVX0 U1096 (.INP(n1031), .ZN(n1107));
   INVX0 U1097 (.INP(n607), .ZN(n1062));
   INVX0 U1098 (.INP(n607), .ZN(n1063));
   INVX0 U1099 (.INP(n623), .ZN(n1038));
   INVX0 U1100 (.INP(n623), .ZN(n1039));
   INVX0 U1101 (.INP(n624), .ZN(n1035));
   INVX0 U1102 (.INP(n624), .ZN(n1036));
   INVX0 U1103 (.INP(n625), .ZN(n1032));
   INVX0 U1104 (.INP(n625), .ZN(n1033));
   INVX0 U1105 (.INP(n626), .ZN(n1029));
   INVX0 U1106 (.INP(n626), .ZN(n1030));
   INVX0 U1107 (.INP(n610), .ZN(n1059));
   INVX0 U1108 (.INP(n610), .ZN(n1060));
   INVX0 U1109 (.INP(n612), .ZN(n1056));
   INVX0 U1110 (.INP(n612), .ZN(n1057));
   INVX0 U1111 (.INP(n613), .ZN(n1053));
   INVX0 U1112 (.INP(n613), .ZN(n1054));
   INVX0 U1113 (.INP(n617), .ZN(n1050));
   INVX0 U1114 (.INP(n617), .ZN(n1051));
   INVX0 U1115 (.INP(n619), .ZN(n1047));
   INVX0 U1116 (.INP(n619), .ZN(n1048));
   INVX0 U1117 (.INP(n620), .ZN(n1044));
   INVX0 U1118 (.INP(n620), .ZN(n1045));
   INVX0 U1119 (.INP(n621), .ZN(n1041));
   INVX0 U1120 (.INP(n621), .ZN(n1042));
   INVX0 U1121 (.INP(n607), .ZN(n1064));
   INVX0 U1122 (.INP(n610), .ZN(n1061));
   INVX0 U1123 (.INP(n612), .ZN(n1058));
   INVX0 U1124 (.INP(n613), .ZN(n1055));
   INVX0 U1125 (.INP(n623), .ZN(n1040));
   INVX0 U1126 (.INP(n624), .ZN(n1037));
   INVX0 U1127 (.INP(n625), .ZN(n1034));
   INVX0 U1128 (.INP(n626), .ZN(n1031));
   INVX0 U1129 (.INP(n617), .ZN(n1052));
   INVX0 U1130 (.INP(n619), .ZN(n1049));
   INVX0 U1131 (.INP(n620), .ZN(n1046));
   INVX0 U1132 (.INP(n621), .ZN(n1043));
   NBUFFX2 U1133 (.INP(n1077), .Z(n1067));
   NBUFFX2 U1134 (.INP(n1077), .Z(n1068));
   NBUFFX2 U1135 (.INP(n1077), .Z(n1069));
   NBUFFX2 U1136 (.INP(n1076), .Z(n1070));
   NBUFFX2 U1137 (.INP(n1076), .Z(n1071));
   NBUFFX2 U1138 (.INP(n1076), .Z(n1072));
   NBUFFX2 U1139 (.INP(n1075), .Z(n1073));
   NBUFFX2 U1140 (.INP(n1075), .Z(n1074));
   NBUFFX2 U1141 (.INP(n1091), .Z(n1081));
   NBUFFX2 U1142 (.INP(n1091), .Z(n1082));
   NBUFFX2 U1143 (.INP(n1091), .Z(n1083));
   NBUFFX2 U1144 (.INP(n1090), .Z(n1084));
   NBUFFX2 U1145 (.INP(n1090), .Z(n1085));
   NBUFFX2 U1146 (.INP(n1090), .Z(n1086));
   NBUFFX2 U1147 (.INP(n1089), .Z(n1087));
   NBUFFX2 U1148 (.INP(n1089), .Z(n1088));
   NBUFFX2 U1149 (.INP(n1105), .Z(n1095));
   NBUFFX2 U1150 (.INP(n1105), .Z(n1096));
   NBUFFX2 U1151 (.INP(n1105), .Z(n1097));
   NBUFFX2 U1152 (.INP(n1104), .Z(n1098));
   NBUFFX2 U1153 (.INP(n1104), .Z(n1099));
   NBUFFX2 U1154 (.INP(n1104), .Z(n1100));
   NBUFFX2 U1155 (.INP(n1103), .Z(n1101));
   NBUFFX2 U1156 (.INP(n1103), .Z(n1102));
   NBUFFX2 U1157 (.INP(n1078), .Z(n1065));
   NBUFFX2 U1158 (.INP(n1078), .Z(n1066));
   NBUFFX2 U1159 (.INP(n1092), .Z(n1079));
   NBUFFX2 U1160 (.INP(n1092), .Z(n1080));
   NBUFFX2 U1161 (.INP(n1106), .Z(n1093));
   NBUFFX2 U1162 (.INP(n1106), .Z(n1094));
   NBUFFX2 U1163 (.INP(n1028), .Z(n1026));
   NBUFFX2 U1164 (.INP(n1078), .Z(n1027));
   NBUFFX2 U1165 (.INP(n1075), .Z(n1028));
   INVX0 U1166 (.INP(n1014), .ZN(n1132));
   INVX0 U1167 (.INP(n1014), .ZN(n1131));
   INVX0 U1168 (.INP(n1016), .ZN(n1137));
   INVX0 U1169 (.INP(n1016), .ZN(n1138));
   INVX0 U1170 (.INP(n1017), .ZN(n1140));
   INVX0 U1171 (.INP(n1017), .ZN(n1141));
   INVX0 U1172 (.INP(n1015), .ZN(n1135));
   INVX0 U1173 (.INP(n1015), .ZN(n1134));
   INVX0 U1174 (.INP(n1014), .ZN(n1133));
   INVX0 U1175 (.INP(n1015), .ZN(n1136));
   INVX0 U1176 (.INP(n1016), .ZN(n1139));
   INVX0 U1177 (.INP(n1017), .ZN(n1142));
   NOR2X0 U1178 (.IN1(n599), .IN2(n588), .QN(n565));
   NOR2X0 U1179 (.IN1(n589), .IN2(n588), .QN(n555));
   NBUFFX2 U1180 (.INP(n1143), .Z(n1077));
   NBUFFX2 U1181 (.INP(n1143), .Z(n1076));
   NBUFFX2 U1182 (.INP(n1143), .Z(n1075));
   NBUFFX2 U1183 (.INP(n1144), .Z(n1091));
   NBUFFX2 U1184 (.INP(n1144), .Z(n1090));
   NBUFFX2 U1185 (.INP(n1144), .Z(n1089));
   NBUFFX2 U1186 (.INP(n1145), .Z(n1105));
   NBUFFX2 U1187 (.INP(n1145), .Z(n1104));
   NBUFFX2 U1188 (.INP(n1145), .Z(n1103));
   NBUFFX2 U1189 (.INP(n1143), .Z(n1078));
   NBUFFX2 U1190 (.INP(n1144), .Z(n1092));
   NBUFFX2 U1191 (.INP(n1145), .Z(n1106));
   NOR2X0 U1192 (.IN1(n1160), .IN2(n1161), .QN(n609));
   INVX0 U1193 (.INP(n616), .ZN(n1153));
   INVX0 U1194 (.INP(n599), .ZN(n1157));
   AO22X1 U1195 (.IN1(n1153), .IN2(write_data[0]), .IN3(core_keylen), .IN4(n616), .Q(n757)
          );
   AO22X1 U1196 (.IN1(n1153), .IN2(write_data[1]), .IN3(core_encdec), .IN4(n616), .Q(n756)
          );
   INVX0 U1197 (.INP(we), .ZN(n1156));
   NOR2X0 U1198 (.IN1(n1160), .IN2(address[0]), .QN(n611));
   NOR2X0 U1199 (.IN1(n1161), .IN2(address[1]), .QN(n598));
   NOR2X0 U1200 (.IN1(address[0]), .IN2(address[1]), .QN(n614));
   NOR2X0 U1201 (.IN1(n627), .IN2(address[2]), .QN(n592));
   INVX0 U1202 (.INP(address[1]), .ZN(n1160));
   INVX0 U1203 (.INP(address[0]), .ZN(n1161));
   NOR2X0 U1204 (.IN1(n1154), .IN2(we), .QN(n606));
   INVX0 U1205 (.INP(n588), .ZN(n1155));
   NAND2X1 U1206 (.IN1(N109), .IN2(N108), .QN(n600));
   AO222X1 U1207 (.IN1(result_reg[2]), .IN2(n1136), .IN3(core_encdec), .IN4(n565), .IN5(
          result_reg[34]), .IN6(n1133), .Q(n568));
   AO222X1 U1208 (.IN1(result_reg[3]), .IN2(n1136), .IN3(core_keylen), .IN4(n565), .IN5(
          result_reg[35]), .IN6(n1133), .Q(n564));
   INVX0 U1209 (.INP(cs), .ZN(n1154));
   INVX0 U1210 (.INP(address[2]), .ZN(n1159));
   NAND2X1 U1211 (.IN1(n596), .IN2(n597), .QN(read_data[0]));
   NAND2X1 U1212 (.IN1(n579), .IN2(n580), .QN(read_data[1]));
   INVX0 U1213 (.INP(address[3]), .ZN(n1158));
   OR2X1 U1214 (.IN1(address[3]), .IN2(address[2]), .Q(n1147));
   AND3X1 U1215 (.IN1(address[4]), .IN2(n1147), .IN3(address[5]), .Q(n1148));
   NOR3X0 U1216 (.IN1(n1148), .IN2(address[7]), .IN3(address[6]), .QN(N109));
   AND2X1 U1217 (.IN1(address[5]), .IN2(address[4]), .Q(n1149));
   OR3X1 U1218 (.IN1(address[7]), .IN2(address[6]), .IN3(n1149), .Q(N108));
   AND2X1 U1219 (.IN1(address[5]), .IN2(address[4]), .Q(n1151));
   OA21X1 U1220 (.IN1(address[3]), .IN2(address[2]), .IN3(address[5]), .Q(n1150));
   NOR4X0 U1221 (.IN1(address[7]), .IN2(address[6]), .IN3(n1151), .IN4(n1150), .QN(N64));
   AND2X1 U1222 (.IN1(address[4]), .IN2(address[3]), .Q(n1152));
   NOR4X0 U1223 (.IN1(address[7]), .IN2(address[6]), .IN3(address[5]), .IN4(n1152), .QN(
          N62));
   aes_DFT_clk_mux_0 occ_snps_pll_controller (.fast_clk(clk), .scan_en(TEST_SE_buf_net1), .
          test_mode(n1560), .reset(pll_reset), .pll_bypass(pll_bypass), .slow_clk(scan_clk)
          , .clk_enable({\clk_ctrl_data[3] , \clk_ctrl_data[2] , \clk_ctrl_data[1] , 
          \clk_ctrl_data[0] }), .clk(n1562));
   aes_DFT_clk_chain_0 snps_clk_chain_0 (.clk(n1562_buf_net1), .se(TEST_SE_buf_net1), .si(
          TEST_SI2), .so(TEST_SO2), .clk_ctrl_data({\clk_ctrl_data[3] , \clk_ctrl_data[2] 
          , \clk_ctrl_data[1] , \clk_ctrl_data[0] }));
   INVX0 U1224 (.INP(SCAN_MODE), .ZN(n1560));
   assign TEST_SE_buf_net0 = TEST_SE;
   assign TEST_SE_buf_net1 = TEST_SE_buf_net0;
   assign n1562_buf_net0 = n1562;
   assign n1562_buf_net1 = n1562_buf_net0;
endmodule

